magic
tech sky130A
magscale 1 2
timestamp 1707921015
<< nwell >>
rect -3160 640 -2740 880
rect -1049 549 -840 870
rect -400 549 -260 870
<< pwell >>
rect -3120 1600 72 5420
<< psubdiff >>
rect -3084 5350 -2988 5384
rect -60 5350 36 5384
rect -3084 5288 -3050 5350
rect -3084 1670 -3050 1732
rect 2 5288 36 5350
rect 2 1670 36 1732
rect -3084 1636 -2988 1670
rect -60 1636 36 1670
<< nsubdiff >>
rect -3060 770 -2960 790
rect -3060 730 -3030 770
rect -2990 730 -2960 770
rect -3060 700 -2960 730
<< psubdiffcont >>
rect -2988 5350 -60 5384
rect -3084 1732 -3050 5288
rect 2 1732 36 5288
rect -2988 1636 -60 1670
<< nsubdiffcont >>
rect -3030 730 -2990 770
<< locali >>
rect -3084 5350 -2988 5384
rect -60 5350 36 5384
rect -3084 5288 -3050 5350
rect -3084 1670 -3050 1732
rect 2 5288 36 5350
rect -1460 1670 -1340 1680
rect 2 1670 36 1732
rect -3084 1636 -2988 1670
rect -60 1636 36 1670
rect -3060 780 -2960 790
rect -3060 730 -3050 780
rect -2980 730 -2960 780
rect -3060 700 -2960 730
<< viali >>
rect -3050 770 -2980 780
rect -3050 730 -3030 770
rect -3030 730 -2990 770
rect -2990 730 -2980 770
rect -120 660 -80 1220
rect -2860 500 -2820 560
rect -830 500 -790 540
rect -2580 430 -2520 470
rect -1140 380 -1080 440
rect -120 -40 -80 120
<< metal1 >>
rect -2940 4820 -2720 5220
rect -2580 4820 -2360 5220
rect -2260 4820 -2040 5220
rect -1920 4820 -1700 5220
rect -1440 4820 -1220 5220
rect -1100 4820 -880 5220
rect -780 4820 -560 5220
rect -440 4820 -220 5220
rect -140 5160 60 5360
rect -140 5000 -20 5160
rect -140 4920 -120 5000
rect -20 4920 -10 5000
rect -2980 3820 -2860 3900
rect -3180 3620 -2860 3820
rect -2980 3480 -2860 3620
rect -2760 3480 -2540 3880
rect -2420 3480 -2200 3880
rect -2100 3480 -1880 3880
rect -1740 3860 -1400 3880
rect -1740 3500 -1620 3860
rect -1540 3500 -1400 3860
rect -1740 3480 -1400 3500
rect -1260 3480 -1040 3880
rect -940 3480 -720 3880
rect -620 3480 -400 3880
rect -300 3440 -220 3520
rect -720 3420 -220 3440
rect -720 3360 -700 3420
rect -620 3360 -220 3420
rect -310 3280 -300 3300
rect -2910 3180 -2900 3280
rect -2800 3200 -1620 3280
rect -1540 3200 -300 3280
rect -2800 3180 -300 3200
rect -180 3180 -170 3300
rect -2890 2660 -2880 3060
rect -2820 2660 -2810 3060
rect -2700 2660 -2520 3040
rect -2360 2660 -2180 3040
rect -2040 2660 -1860 3040
rect -1700 2920 -940 2940
rect -1700 2700 -1040 2920
rect -940 2700 -930 2920
rect -2860 1820 -2680 2200
rect -2520 1820 -2340 2200
rect -2200 1820 -2020 2200
rect -1860 2120 -1680 2200
rect 6280 2160 6500 2180
rect 6280 2120 6300 2160
rect -1860 2000 -1660 2120
rect -1050 2020 -1040 2120
rect -920 2020 -300 2120
rect -1040 2000 -300 2020
rect -220 2000 6300 2120
rect -1860 1820 -1680 2000
rect 6280 1980 6300 2000
rect 6480 2120 6500 2160
rect 6480 2000 6950 2120
rect 6480 1980 6500 2000
rect 6280 1960 6500 1980
rect -310 1280 -300 1340
rect -240 1320 -230 1340
rect -240 1280 -220 1320
rect -3180 1190 -2980 1240
rect -3180 1080 -580 1190
rect -510 1080 -500 1190
rect -3180 1040 -2980 1080
rect -3180 880 -2980 940
rect -3180 780 -2840 880
rect -3180 740 -3050 780
rect -3060 730 -3050 740
rect -2980 730 -2960 780
rect -3060 700 -2960 730
rect -410 660 -400 1240
rect -340 660 -300 1240
rect -126 1220 -74 1232
rect -220 660 -120 1220
rect -80 1200 -40 1220
rect -40 1120 -30 1200
rect -80 1080 -40 1120
rect -40 1000 -30 1080
rect -80 940 -40 1000
rect -40 860 -30 940
rect -80 800 -40 860
rect -40 720 -30 800
rect -80 660 -40 720
rect -126 648 -74 660
rect -3180 560 -2980 600
rect -2866 560 -2814 572
rect -3180 500 -2860 560
rect -2820 500 -2814 560
rect -3180 400 -2980 500
rect -2866 488 -2814 500
rect -842 540 -778 546
rect -590 540 -580 560
rect -842 500 -830 540
rect -790 500 -580 540
rect -842 494 -778 500
rect -590 480 -580 500
rect -500 480 -490 560
rect -300 540 -280 580
rect -290 520 -280 540
rect -220 520 -210 580
rect -2600 410 -2590 480
rect -2510 410 -2500 480
rect -2150 420 -2140 480
rect -2080 420 -2070 480
rect -1152 440 -1068 446
rect -1152 380 -1140 440
rect -1080 380 -700 440
rect -620 380 -610 440
rect -1152 374 -1068 380
rect -2870 240 -2860 320
rect -2780 240 -2770 320
rect -290 240 -280 260
rect -300 200 -280 240
rect -220 200 -210 260
rect -2590 140 -2580 200
rect -2520 190 -350 200
rect -2520 140 -420 190
rect -430 130 -420 140
rect -360 140 -350 190
rect -360 130 -300 140
rect -3180 -20 -2980 40
rect -3180 -80 -2140 -20
rect -2080 -80 -2070 -20
rect -410 -40 -300 130
rect -220 120 -20 140
rect -220 100 -120 120
rect -80 100 -20 120
rect -220 -40 -160 100
rect -60 -40 -20 100
rect -140 -60 -20 -40
rect -3180 -160 -2980 -80
rect -300 -120 -220 -80
rect -1760 -360 -1560 -320
rect -2900 -500 -2880 -360
rect -2780 -380 -60 -360
rect -2780 -500 -160 -380
rect -60 -500 -50 -380
rect -2900 -520 -60 -500
<< via1 >>
rect -120 4920 -20 5000
rect -1620 3500 -1540 3860
rect -700 3360 -620 3420
rect -2900 3180 -2800 3280
rect -1620 3200 -1540 3280
rect -300 3180 -180 3300
rect -2880 2660 -2820 3060
rect -1040 2700 -940 2920
rect -1040 2020 -920 2120
rect -300 2000 -220 2120
rect 6300 1980 6480 2160
rect -300 1280 -240 1340
rect -580 1080 -510 1190
rect -400 660 -340 1240
rect -120 1120 -80 1200
rect -80 1120 -40 1200
rect -120 1000 -80 1080
rect -80 1000 -40 1080
rect -120 860 -80 940
rect -80 860 -40 940
rect -120 720 -80 800
rect -80 720 -40 800
rect -580 480 -500 560
rect -280 520 -220 580
rect -2590 470 -2510 480
rect -2590 430 -2580 470
rect -2580 430 -2520 470
rect -2520 430 -2510 470
rect -2590 410 -2510 430
rect -2140 420 -2080 480
rect -700 380 -620 440
rect -2860 240 -2780 320
rect -280 200 -220 260
rect -2580 140 -2520 200
rect -420 130 -360 190
rect -2140 -80 -2080 -20
rect -160 -40 -120 100
rect -120 -40 -80 100
rect -80 -40 -60 100
rect -2880 -500 -2780 -360
rect -160 -500 -60 -380
<< metal2 >>
rect -120 5000 -20 5010
rect -140 4920 -120 5000
rect -1620 3860 -1520 3880
rect -1540 3500 -1520 3860
rect -2900 3280 -2800 3290
rect -2900 3060 -2800 3180
rect -1620 3280 -1520 3500
rect -1540 3200 -1520 3280
rect -1620 3160 -1520 3200
rect -700 3420 -620 3430
rect -2900 2660 -2880 3060
rect -2820 2660 -2800 3060
rect -2900 2640 -2800 2660
rect -1040 2920 -920 2960
rect -940 2700 -920 2920
rect -1040 2120 -920 2700
rect -1040 2000 -920 2020
rect -2590 480 -2510 490
rect -2590 400 -2510 410
rect -2140 480 -2080 490
rect -2860 320 -2780 330
rect -2880 240 -2860 320
rect -2880 -360 -2780 240
rect -2580 210 -2540 400
rect -2580 200 -2520 210
rect -2580 130 -2520 140
rect -2140 -20 -2080 420
rect -700 440 -620 3360
rect -300 3300 -180 3310
rect -300 3170 -180 3180
rect -300 2120 -220 2130
rect -300 1340 -220 2000
rect -240 1280 -220 1340
rect -300 1270 -240 1280
rect -400 1240 -340 1250
rect -580 1190 -510 1200
rect -580 570 -510 1080
rect -140 1200 -20 4920
rect 6280 2160 6500 2180
rect 6280 1980 6300 2160
rect 6480 1980 6500 2160
rect 6280 1960 6500 1980
rect -140 1120 -120 1200
rect -40 1120 -20 1200
rect -140 1080 -20 1120
rect -140 1000 -120 1080
rect -40 1000 -20 1080
rect -140 940 -20 1000
rect -140 860 -120 940
rect -40 860 -20 940
rect -140 800 -20 860
rect -140 720 -120 800
rect -40 720 -20 800
rect -140 660 -20 720
rect -580 560 -500 570
rect -580 470 -500 480
rect -700 370 -620 380
rect -400 200 -340 660
rect -420 190 -340 200
rect -280 580 -220 590
rect -280 260 -220 520
rect -280 190 -220 200
rect -360 130 -340 190
rect -420 120 -340 130
rect -400 -40 -340 120
rect -160 100 -60 280
rect -2140 -90 -2080 -80
rect -2880 -510 -2780 -500
rect -160 -380 -60 -40
rect -160 -510 -60 -500
<< via2 >>
rect -300 3180 -180 3300
rect 6300 1980 6480 2160
rect -160 -480 -60 -380
<< metal3 >>
rect -320 3300 -160 3320
rect -320 3180 -300 3300
rect -180 3180 -160 3300
rect -320 3160 -160 3180
rect 6280 2160 6500 2180
rect 6280 1980 6300 2160
rect 6480 1980 6500 2160
rect 6280 1960 6500 1980
rect -200 -380 7100 -360
rect -200 -480 -160 -380
rect -60 -480 7100 -380
rect -200 -520 7100 -480
<< via3 >>
rect -300 3180 -180 3300
rect 6300 1980 6480 2160
<< metal4 >>
rect -540 3300 500 3320
rect -540 3180 -300 3300
rect -180 3180 500 3300
rect -540 2880 500 3180
rect 6440 2180 7300 2280
rect 6280 2160 7300 2180
rect 6280 1980 6300 2160
rect 6480 1980 7300 2160
rect 6280 1960 7300 1980
rect 6440 1840 7300 1960
<< comment >>
rect 220 -500 240 -480
rect 6600 -500 6620 -480
rect 6120 -520 6140 -500
use sky130_fd_pr__cap_mim_m3_1_A4KLY5  sky130_fd_pr__cap_mim_m3_1_A4KLY5_0
timestamp 1707920920
transform 0 1 9380 -1 0 2426
box -2906 -2760 2906 2760
use sky130_fd_pr__cap_mim_m3_1_A4KLY5  sky130_fd_pr__cap_mim_m3_1_A4KLY5_1
timestamp 1707920920
transform 0 1 3000 -1 0 2426
box -2906 -2760 2906 2760
use sky130_fd_pr__nfet_01v8_648S5X  sky130_fd_pr__nfet_01v8_648S5X_0
timestamp 1700078798
transform 1 0 -255 0 1 54
box -211 -310 211 310
use sky130_fd_pr__res_xhigh_po_0p35_QABHPF  sky130_fd_pr__res_xhigh_po_0p35_QABHPF_0
timestamp 1701394307
transform 1 0 -2264 0 1 2432
box -616 -632 616 632
use sky130_fd_pr__res_xhigh_po_0p35_XMXTTL  sky130_fd_pr__res_xhigh_po_0p35_XMXTTL_1
timestamp 1700079212
transform 1 0 -2314 0 1 4350
box -616 -882 616 882
use sky130_fd_pr__res_xhigh_po_0p35_XMXTTL  sky130_fd_pr__res_xhigh_po_0p35_XMXTTL_2
timestamp 1700079212
transform 1 0 -840 0 1 4350
box -616 -882 616 882
use sky130_fd_sc_hd__dfrbp_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 -2882 0 1 288
box -38 -48 2154 592
use sky130_fd_pr__pfet_01v8_XGSNAL  XP1
timestamp 1700078798
transform 1 0 -255 0 1 933
box -211 -519 211 519
<< labels >>
flabel metal1 -3180 740 -2980 940 0 FreeSans 1600 0 0 0 vpwr
port 2 nsew
flabel metal1 -3180 400 -2980 600 0 FreeSans 1600 0 0 0 clk
port 3 nsew
flabel metal1 -3180 -160 -2980 40 0 FreeSans 1600 0 0 0 reset_b_dff
port 4 nsew
flabel metal1 -1760 -520 -1560 -320 0 FreeSans 1600 0 0 0 gnd
port 6 nsew
flabel metal1 -140 5160 60 5360 0 FreeSans 1600 0 0 0 vd
port 8 nsew
flabel metal1 -1400 3220 -1340 3240 0 FreeSans 800 0 0 0 in_int
flabel metal1 -1340 2820 -1280 2840 0 FreeSans 800 0 0 0 in_comp
flabel metal1 -3180 1040 -2980 1240 0 FreeSans 1600 0 0 0 out
port 1 nsew
flabel metal1 -3180 3620 -2980 3820 0 FreeSans 1600 0 0 0 in
port 9 nsew
<< end >>
