* NGSPICE file created from tt_um_hugodiasg_temp-sensor_clock-divider.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_FRXWNM a_n100_n297# a_100_n200# w_n194_n300# a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n194_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_FVXEPM a_n100_n297# a_100_n200# w_n194_n300# a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n194_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_FVTXNM a_29_n297# a_n287_n200# a_n229_n297# a_229_n200#
+ a_n29_n200# w_n323_n300#
X0 a_229_n200# a_29_n297# a_n29_n200# w_n323_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X1 a_n29_n200# a_n229_n297# a_n287_n200# w_n323_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_3HGYVM a_n100_n297# a_100_n200# w_n194_n300# a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n194_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_SKTYVM a_n500_n297# a_500_n200# w_n594_n300# a_n558_n200#
X0 a_500_n200# a_n500_n297# a_n558_n200# w_n594_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=5
.ends

.subckt sky130_fd_pr__nfet_01v8_9VJR3B a_100_527# a_n158_n727# a_100_n309# a_n100_21#
+ a_n158_n309# a_100_109# a_n158_527# a_n100_n815# a_n100_439# a_n158_109# a_100_n727#
+ a_n100_n397# VSUBS
X0 a_100_n309# a_n100_n397# a_n158_n309# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_527# a_n100_439# a_n158_527# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_n727# a_n100_n815# a_n158_n727# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_109# a_n100_21# a_n158_109# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_YAWWFM a_29_n297# a_n287_n200# w_n581_n300# a_n229_n297#
+ a_287_n297# a_229_n200# a_n545_n200# a_n487_n297# a_487_n200# a_n29_n200#
X0 a_229_n200# a_29_n297# a_n29_n200# w_n581_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_n29_n200# a_n229_n297# a_n287_n200# w_n581_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_n287_n200# a_n487_n297# a_n545_n200# w_n581_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X3 a_487_n200# a_287_n297# a_229_n200# w_n581_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_YAEUFM a_29_n297# a_n287_n200# a_n1061_n200# a_n745_n297#
+ a_745_n200# a_803_n297# a_n229_n297# a_n1003_n297# a_287_n297# a_229_n200# a_n545_n200#
+ a_1003_n200# a_n487_n297# a_487_n200# a_n29_n200# a_545_n297# a_n803_n200# w_n1097_n300#
X0 a_229_n200# a_29_n297# a_n29_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_n29_n200# a_n229_n297# a_n287_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_n545_n200# a_n745_n297# a_n803_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_n287_n200# a_n487_n297# a_n545_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_n803_n200# a_n1003_n297# a_n1061_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X5 a_1003_n200# a_803_n297# a_745_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X6 a_745_n200# a_545_n297# a_487_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_487_n200# a_287_n297# a_229_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sensor vd vts vtd gnd
Xsky130_fd_pr__pfet_01v8_FRXWNM_0 vd vd vd vd sky130_fd_pr__pfet_01v8_FRXWNM
Xsky130_fd_pr__pfet_01v8_FRXWNM_1 vd vd vd vd sky130_fd_pr__pfet_01v8_FRXWNM
Xsky130_fd_pr__pfet_01v8_FVXEPM_0 c c vd c sky130_fd_pr__pfet_01v8_FVXEPM
Xsky130_fd_pr__pfet_01v8_FRXWNM_2 vd vd vd vd sky130_fd_pr__pfet_01v8_FRXWNM
Xsky130_fd_pr__pfet_01v8_FRXWNM_3 vts vts vts vts sky130_fd_pr__pfet_01v8_FRXWNM
Xsky130_fd_pr__pfet_01v8_FRXWNM_4 vts vts vts vts sky130_fd_pr__pfet_01v8_FRXWNM
XXP1 a a a a vd vd sky130_fd_pr__pfet_01v8_FVTXNM
XXP3 vtd d vd vd sky130_fd_pr__pfet_01v8_3HGYVM
XXP4 vtd vd vd vts sky130_fd_pr__pfet_01v8_SKTYVM
Xsky130_fd_pr__nfet_01v8_9VJR3B_0 gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd
+ gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_2 a gnd a b gnd a gnd b b gnd a b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_1 gnd a gnd b a gnd a b b a gnd b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_3 gnd vtd gnd b vtd gnd vtd b b vtd gnd b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_4 vtd gnd vtd b gnd vtd gnd b b gnd vtd b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_5 gnd b gnd b b gnd b b b b gnd b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_6 gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd
+ gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__pfet_01v8_YAWWFM_1 vtd b vd vtd vtd b c vtd c c sky130_fd_pr__pfet_01v8_YAWWFM
Xsky130_fd_pr__pfet_01v8_YAWWFM_0 a d vd a a d c a c c sky130_fd_pr__pfet_01v8_YAWWFM
Xsky130_fd_pr__nfet_01v8_9VJR3B_7 b gnd b b gnd b gnd b b gnd b b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__pfet_01v8_YAEUFM_0 vtd vts vtd vtd vts vtd vtd vtd vtd vts vtd vtd
+ vtd vtd vtd vtd vts vts sky130_fd_pr__pfet_01v8_YAEUFM
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.106 ps=0.975 w=0.65 l=0.15
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.162 ps=1.33 w=1 l=0.15
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0991 ps=0.955 w=0.65 l=0.15
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.28 ps=1.62 w=1 l=0.15
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0619 ps=0.715 w=0.42 l=0.15
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0746 pd=0.775 as=0.109 ps=1.36 w=0.42 l=0.15
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.62 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.175 ps=1.26 w=0.65 l=0.15
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0746 ps=0.775 w=0.42 l=0.15
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.136 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258 ps=1.45 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.1 as=0.111 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258 pd=1.45 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.272 ps=2.56 w=1 l=0.15
X15 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X17 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X19 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X24 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.257 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X30 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X38 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.185 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
X0 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X36 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_33_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.182 ps=1.86 w=0.65 l=0.15
X4 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X11 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B1_N a_33_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X20 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.162 pd=1.15 as=0.111 ps=0.99 w=0.65 l=0.15
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.162 ps=1.15 w=0.65 l=0.15
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.123 ps=1.03 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.198 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.393 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.393 ps=1.78 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.146 ps=1.34 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.209 pd=1.35 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.209 ps=1.35 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0662 pd=0.735 as=0.0986 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0986 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.266 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.102 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.111 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.119 ps=1.01 w=0.65 l=0.15
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.62 as=0.26 ps=2.52 w=1 l=0.15
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203 pd=1.27 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.312 ps=1.62 w=1 l=0.15
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.137 ps=1.07 w=0.65 l=0.15
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203 ps=1.27 w=0.65 l=0.15
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.21 ps=1.42 w=1 l=0.15
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.138 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.1 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_82_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 a_646_47# B2 a_82_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_574_369# a_313_47# a_82_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0976 pd=0.945 as=0.166 ps=1.8 w=0.64 l=0.15
X3 a_574_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4 VGND a_82_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR B2 a_574_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0976 ps=0.945 w=0.64 l=0.15
X6 X a_82_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X7 X a_82_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8 a_313_47# A2_N a_313_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.0672 ps=0.85 w=0.64 l=0.15
X9 a_313_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 a_313_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.186 ps=1.43 w=0.64 l=0.15
X11 VGND A2_N a_313_47# VNB sky130_fd_pr__nfet_01v8 ad=0.142 pd=1.1 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_82_21# a_313_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.142 ps=1.1 w=0.42 l=0.15
X13 VGND B1 a_646_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.183 ps=1.24 w=0.65 l=0.15
X1 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_479_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X4 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 Y a_61_47# a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_61_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X8 VGND A2 a_637_47# VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_61_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A1 a_479_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0683 ps=0.86 w=0.65 l=0.15
X11 VGND B1_N a_61_47# VNB sky130_fd_pr__nfet_01v8 ad=0.183 pd=1.24 as=0.126 ps=1.44 w=0.42 l=0.15
X12 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X13 a_637_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt clock_divider clk_in clk_out nrst scale[0] scale[1] scale[2] scale[3] scale[4]
+ scale[5] scale[6] scale[7] VPWR VGND
XFILLER_0_17_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0985_ count\[27\] _0486_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_19_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0770_ _0139_ _0293_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__nand2_1
X_0968_ count\[21\] _0474_ _0447_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__o21ai_1
X_0899_ _0427_ _0429_ _0063_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0822_ net16 _0338_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__nor2_1
X_0753_ _0288_ _0289_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0684_ _0207_ _0210_ _0224_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1021_ net22 _0018_ VGND VGND VPWR VPWR true_scale\[23\] sky130_fd_sc_hd__dfxtp_1
X_0805_ net8 net10 net9 VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a21oi_1
X_0598_ _0141_ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__xor2_2
X_0736_ _0271_ _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__xnor2_2
X_0667_ _0208_ _0111_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0521_ net4 _0070_ _0071_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__o21a_1
X_1004_ net19 _0001_ VGND VGND VPWR VPWR true_scale\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0719_ _0241_ _0242_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_33_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0504_ true_scale\[15\] true_scale\[16\] true_scale\[17\] _0057_ VGND VGND VPWR VPWR
+ _0058_ sky130_fd_sc_hd__or4_2
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0984_ _0488_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0967_ count\[19\] count\[20\] count\[21\] _0471_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__and4_1
X_0898_ count\[26\] count\[27\] _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0752_ _0163_ _0287_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__or2_1
X_0821_ _0068_ _0351_ _0352_ _0353_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0683_ _0209_ _0096_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__and2b_1
X_1020_ net22 _0017_ VGND VGND VPWR VPWR true_scale\[22\] sky130_fd_sc_hd__dfxtp_1
X_0804_ net8 net9 net10 VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__and3_1
X_0735_ _0123_ _0253_ _0272_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__o21a_1
X_0666_ _0075_ _0080_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__nand2_1
X_0597_ net4 _0124_ _0092_ _0125_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0520_ net4 net5 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ net19 _0000_ VGND VGND VPWR VPWR true_scale\[5\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0718_ _0139_ _0256_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__xnor2_1
X_0649_ _0190_ _0191_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0503_ true_scale\[12\] true_scale\[13\] true_scale\[14\] _0056_ VGND VGND VPWR VPWR
+ _0057_ sky130_fd_sc_hd__or4_2
XFILLER_0_17_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0983_ _0486_ _0487_ _0432_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__and3b_1
X_0897_ count\[28\] count\[29\] count\[30\] count\[31\] VGND VGND VPWR VPWR _0428_
+ sky130_fd_sc_hd__or4_1
X_0966_ _0476_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
X_0751_ _0163_ _0287_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0820_ true_scale\[25\] net16 VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__and2_1
X_0682_ _0107_ _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0949_ count\[13\] count\[14\] count\[15\] _0459_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__and4_2
XFILLER_0_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0734_ _0127_ _0252_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__nand2_1
X_0803_ _0331_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__inv_2
X_0665_ _0205_ _0206_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__nor2_1
X_0596_ _0072_ _0140_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__xor2_2
XFILLER_0_30_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1002_ _0068_ _0500_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__nor2_1
X_0648_ _0168_ _0170_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0717_ _0254_ _0255_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__xnor2_2
X_0579_ _0066_ _0124_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0502_ true_scale\[9\] true_scale\[10\] true_scale\[11\] _0055_ VGND VGND VPWR VPWR
+ _0056_ sky130_fd_sc_hd__or4_2
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0982_ count\[24\] count\[25\] _0480_ count\[26\] VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0896_ _0425_ _0426_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__nand2_1
X_0965_ _0474_ _0475_ _0437_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__and3b_1
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0750_ _0285_ _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0681_ _0095_ _0220_ _0221_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a21bo_1
X_0948_ _0464_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0879_ true_scale\[21\] _0059_ true_scale\[22\] VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0802_ _0068_ _0334_ _0335_ _0336_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a31o_1
X_0733_ _0146_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__xnor2_2
X_0664_ net10 _0089_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__nor2_1
X_0595_ net7 net13 VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__xor2_4
XFILLER_0_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1001_ signal_clk_out _0431_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__xor2_1
X_0647_ _0185_ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__xnor2_2
X_0716_ _0113_ _0146_ _0130_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__a21oi_2
X_0578_ net14 net5 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0501_ true_scale\[5\] true_scale\[6\] true_scale\[7\] true_scale\[8\] VGND VGND
+ VPWR VPWR _0055_ sky130_fd_sc_hd__or4_2
XFILLER_0_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0981_ count\[25\] count\[26\] _0483_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0964_ count\[19\] _0471_ count\[20\] VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__a21o_1
X_0895_ count\[28\] count\[29\] VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0680_ _0111_ _0094_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__nand2_1
X_0947_ _0462_ _0463_ _0437_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__and3b_1
XFILLER_0_27_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0878_ count\[20\] _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0801_ true_scale\[23\] net16 VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__and2_1
X_0594_ _0138_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__buf_4
X_0732_ _0268_ _0269_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__xnor2_2
X_0663_ net6 net7 net10 VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1000_ count\[31\] _0496_ _0499_ _0447_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__o211a_1
X_0715_ _0146_ _0253_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__xnor2_2
X_0646_ _0187_ _0188_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0577_ net10 net12 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__xnor2_4
XPHY_EDGE_ROW_11_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_75 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0629_ _0141_ _0142_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__nand2_1
X_0980_ count\[25\] _0483_ _0485_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0894_ count\[26\] count\[27\] count\[30\] count\[31\] VGND VGND VPWR VPWR _0425_
+ sky130_fd_sc_hd__and4_1
X_0963_ count\[19\] count\[20\] _0471_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0946_ count\[13\] _0459_ count\[14\] VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__a21o_1
X_0877_ true_scale\[21\] _0059_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_41_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0800_ _0333_ _0322_ _0323_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__or3_1
X_0731_ _0111_ _0251_ _0080_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__o21a_1
X_0662_ _0145_ _0182_ _0183_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__o21bai_4
X_0593_ net10 _0107_ _0122_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__a21bo_1
X_0929_ _0450_ _0451_ _0437_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__and3b_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0645_ _0082_ _0083_ _0186_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__o21ai_1
X_0714_ _0127_ _0252_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__xnor2_2
X_0576_ net9 _0106_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0628_ _0170_ _0171_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_87 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0559_ net13 _0081_ _0089_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__a21o_2
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0962_ count\[19\] _0471_ _0473_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__a21oi_1
X_0893_ count\[25\] _0423_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0945_ count\[13\] count\[14\] _0459_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__and3_1
X_0876_ count\[19\] _0406_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0661_ _0181_ _0192_ _0202_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0730_ net5 _0140_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__xnor2_2
X_0592_ _0068_ _0135_ _0136_ _0137_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a31o_1
X_0928_ count\[7\] _0446_ count\[8\] VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__a21o_1
X_0859_ _0388_ _0389_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0713_ _0092_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__xnor2_2
X_0644_ _0082_ _0083_ _0186_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__nor3_1
X_0575_ net15 _0119_ _0120_ _0121_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__o31ai_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0627_ _0168_ _0169_ _0163_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0558_ _0095_ _0096_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0961_ count\[19\] _0471_ _0433_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0892_ true_scale\[26\] _0062_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0944_ count\[13\] _0459_ _0461_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ _0059_ _0405_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__nand2_1
X_0660_ _0191_ _0190_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__and2b_1
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0591_ true_scale\[12\] net15 VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ count\[7\] count\[8\] _0446_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0858_ true_scale\[15\] _0057_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__and2_1
X_0789_ _0312_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0574_ true_scale\[11\] net15 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__nand2_1
X_0712_ _0250_ _0093_ _0079_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__or3_2
X_0643_ _0075_ _0165_ _0079_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__a21oi_1
X_1057_ net23 _0054_ VGND VGND VPWR VPWR signal_clk_out sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_15_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0626_ _0163_ _0168_ _0169_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0557_ true_scale\[10\] net15 _0104_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0609_ _0150_ _0153_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__xnor2_1
X_0960_ _0471_ _0472_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0891_ count\[24\] _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_18_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0943_ count\[13\] _0459_ _0433_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__o21ai_1
X_0874_ true_scale\[18\] true_scale\[19\] _0058_ true_scale\[20\] VGND VGND VPWR VPWR
+ _0405_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0590_ _0133_ _0134_ _0103_ _0123_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0926_ count\[7\] _0446_ _0449_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0857_ true_scale\[15\] _0057_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__nor2_1
X_0788_ _0318_ _0314_ _0315_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0711_ net4 net3 VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__nor2_1
X_0642_ _0145_ _0184_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_20_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0573_ _0103_ _0118_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__nor2_1
X_1056_ net20 _0053_ VGND VGND VPWR VPWR count\[31\] sky130_fd_sc_hd__dfxtp_1
X_0909_ count\[0\] count\[1\] count\[2\] VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0625_ _0166_ _0167_ _0079_ _0164_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__a211oi_1
X_0556_ _0090_ _0102_ _0103_ _0068_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__o211a_1
X_1039_ net18 _0036_ VGND VGND VPWR VPWR count\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0608_ _0122_ _0151_ _0152_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__o21a_1
X_0539_ _0084_ _0085_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ _0062_ _0420_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0942_ _0459_ _0460_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__nor2_1
X_0873_ _0394_ _0397_ _0401_ _0403_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0925_ count\[7\] _0446_ _0433_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__o21ai_1
X_0856_ count\[13\] _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0787_ _0299_ _0302_ _0316_ _0317_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0641_ _0182_ _0183_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__nor2_2
X_0710_ _0249_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
X_0572_ _0103_ _0118_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__and2_1
X_1055_ net20 _0052_ VGND VGND VPWR VPWR count\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0908_ _0432_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__buf_2
X_0839_ _0368_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0624_ _0079_ _0164_ _0166_ _0167_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__o211a_1
X_0555_ _0090_ _0095_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__nand2_1
X_1038_ net18 _0035_ VGND VGND VPWR VPWR count\[13\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0538_ net6 _0079_ _0086_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__a21o_1
X_0607_ _0131_ _0129_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout20 net21 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0941_ count\[12\] _0456_ _0447_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__o21ai_1
X_0872_ count\[18\] _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0924_ _0446_ _0448_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0855_ _0057_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nand2_1
X_0786_ _0321_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0640_ net6 net13 net9 VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__and3_1
X_0571_ _0100_ _0117_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__xnor2_1
X_1054_ net20 _0051_ VGND VGND VPWR VPWR count\[29\] sky130_fd_sc_hd__dfxtp_1
X_0907_ count\[0\] count\[1\] count\[2\] VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0838_ true_scale\[9\] _0055_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__and2_1
X_0769_ _0305_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0623_ _0075_ _0080_ _0165_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0554_ _0100_ _0101_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__nor2_1
X_1037_ net18 _0034_ VGND VGND VPWR VPWR count\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0537_ _0084_ _0085_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__nand2_1
X_0606_ _0129_ _0131_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__and2b_1
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout21 net23 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0940_ count\[10\] count\[11\] count\[12\] _0453_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__and4_2
XFILLER_0_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0871_ true_scale\[19\] _0398_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0923_ count\[6\] _0443_ _0447_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__o21ai_1
X_0854_ true_scale\[12\] true_scale\[13\] _0056_ true_scale\[14\] VGND VGND VPWR VPWR
+ _0385_ sky130_fd_sc_hd__o31ai_1
X_0785_ true_scale\[22\] _0320_ _0067_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_7_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0570_ _0115_ _0116_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__and2b_1
X_1053_ net20 _0050_ VGND VGND VPWR VPWR count\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0906_ count\[0\] count\[1\] _0435_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__o21a_1
X_0837_ true_scale\[9\] _0055_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__nor2_1
X_0768_ true_scale\[21\] _0304_ _0067_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
X_0699_ _0223_ _0225_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0553_ _0098_ _0099_ _0086_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__o21a_1
X_0622_ _0075_ _0080_ _0165_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__a21o_1
X_1036_ net18 _0033_ VGND VGND VPWR VPWR count\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0605_ _0139_ _0149_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__xnor2_2
X_0536_ net6 _0075_ _0079_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ net22 _0016_ VGND VGND VPWR VPWR true_scale\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0519_ net14 net5 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__xor2_1
Xfanout22 net23 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ count\[17\] _0400_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__xnor2_1
X_0999_ count\[30\] count\[31\] _0426_ _0489_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__nand4_1
XFILLER_0_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0922_ _0432_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__buf_2
X_0853_ _0374_ _0377_ _0381_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__or4_1
X_0784_ _0316_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__xnor2_1
Xinput1 clk_in VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1052_ net20 _0049_ VGND VGND VPWR VPWR count\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0905_ count\[0\] count\[1\] _0433_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__a21boi_1
X_0836_ _0365_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__or2_1
X_0767_ _0297_ _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__xnor2_1
X_0698_ _0238_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
X_0621_ net6 net13 VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__xor2_4
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0552_ _0086_ _0098_ _0099_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__nor3_1
X_1035_ net18 _0032_ VGND VGND VPWR VPWR count\[10\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_10_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0819_ _0348_ _0350_ _0347_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0604_ _0144_ _0148_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__xor2_2
X_0535_ _0082_ _0083_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1018_ net22 _0015_ VGND VGND VPWR VPWR true_scale\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0518_ _0069_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__clkbuf_1
Xfanout23 net1 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_41_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0998_ _0498_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
X_0921_ count\[4\] count\[5\] count\[6\] _0355_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__and4_2
XFILLER_0_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0852_ count\[12\] _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0783_ _0317_ _0303_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 nrst VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_40_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1051_ net20 _0048_ VGND VGND VPWR VPWR count\[26\] sky130_fd_sc_hd__dfxtp_1
X_0904_ _0434_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0835_ _0055_ _0364_ count\[7\] VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__a21oi_1
X_0697_ true_scale\[17\] _0237_ _0067_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux2_1
X_0766_ _0299_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0551_ _0089_ _0097_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__nor2_1
X_0620_ net4 _0070_ _0140_ _0071_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__o211a_1
X_1034_ net17 _0031_ VGND VGND VPWR VPWR count\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0749_ net5 _0140_ _0165_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__nand3_1
X_0818_ _0347_ _0348_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0534_ _0075_ _0080_ _0081_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__a21oi_1
X_0603_ _0146_ _0128_ _0147_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__a21o_1
X_1017_ net22 _0014_ VGND VGND VPWR VPWR true_scale\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0517_ true_scale\[6\] _0066_ _0068_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_1
Xfanout13 net8 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_8
XFILLER_0_35_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0997_ _0496_ _0437_ _0497_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__and3b_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0920_ _0445_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
X_0851_ true_scale\[13\] _0378_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0782_ _0294_ _0296_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 scale[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ net21 _0047_ VGND VGND VPWR VPWR count\[25\] sky130_fd_sc_hd__dfxtp_1
X_0903_ count\[0\] _0433_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__and2b_1
X_0834_ count\[7\] _0055_ _0364_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__and3_1
X_0696_ _0230_ _0236_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__xnor2_1
X_0765_ _0279_ _0300_ _0298_ _0263_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0550_ _0089_ _0097_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__and2_1
X_1033_ net17 _0030_ VGND VGND VPWR VPWR count\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0817_ _0322_ _0323_ _0349_ _0333_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__o211a_1
X_0748_ net5 _0140_ _0165_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__a21o_1
X_0679_ _0208_ _0111_ _0080_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0533_ _0075_ _0080_ _0081_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0602_ _0126_ _0127_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1016_ net22 _0013_ VGND VGND VPWR VPWR true_scale\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0516_ _0067_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout14 net3 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0996_ count\[27\] _0426_ _0486_ count\[30\] VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ count\[11\] _0380_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__xnor2_1
X_0781_ _0297_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__inv_2
Xinput4 scale[1] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0979_ count\[25\] _0483_ _0433_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_27_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0902_ _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__buf_2
X_0833_ true_scale\[8\] _0357_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__nand2_1
X_0695_ _0231_ net11 _0234_ _0235_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a211o_1
X_0764_ _0275_ _0277_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1032_ net17 _0029_ VGND VGND VPWR VPWR count\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0747_ _0123_ _0270_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__nor2_1
X_0816_ _0341_ _0342_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__nor2_1
X_0678_ _0219_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
X_0601_ _0145_ net12 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__xnor2_4
X_0532_ net6 net7 VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__xor2_4
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ net22 _0012_ VGND VGND VPWR VPWR true_scale\[17\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_14_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0515_ net16 VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__inv_2
Xfanout15 net2 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XFILLER_0_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ count\[30\] _0426_ _0489_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__and3_1
X_0780_ _0314_ _0315_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__and2b_1
Xinput5 scale[2] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0978_ _0483_ _0484_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_2_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0832_ _0356_ _0359_ _0360_ _0362_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__or4b_1
X_0901_ net16 _0431_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__and2_1
X_0763_ _0275_ _0277_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__nand2_1
X_0694_ _0198_ _0196_ _0197_ _0215_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__nor4_1
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap12 _0107_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_4
X_1031_ net17 _0028_ VGND VGND VPWR VPWR count\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0815_ _0331_ _0342_ _0341_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__o21ba_1
X_0746_ _0268_ _0269_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__nor2_1
X_0677_ true_scale\[16\] _0218_ _0067_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0600_ net10 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__inv_4
X_0531_ net4 net14 net5 VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__nand3_2
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ net22 _0011_ VGND VGND VPWR VPWR true_scale\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0729_ _0068_ _0265_ _0266_ _0267_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_31_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0514_ net4 net14 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__xor2_1
Xfanout16 net2 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
XFILLER_0_36_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0994_ _0494_ _0492_ _0495_ _0447_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 scale[3] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0977_ count\[24\] _0480_ _0447_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0419_ _0422_ _0424_ _0430_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0831_ count\[4\] true_scale\[5\] _0361_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__mux2_1
X_0762_ _0235_ _0234_ net11 _0261_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__o311a_1
X_0693_ _0203_ _0214_ _0233_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1030_ net17 _0027_ VGND VGND VPWR VPWR count\[5\] sky130_fd_sc_hd__dfxtp_1
X_0814_ _0145_ _0338_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__nor2_1
X_0676_ _0215_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__xnor2_1
X_0745_ _0282_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0530_ _0078_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1013_ net1 _0010_ VGND VGND VPWR VPWR true_scale\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0659_ _0201_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
X_0728_ true_scale\[19\] net16 VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__and2_1
X_0513_ _0065_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
Xfanout17 net19 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
X_0993_ _0494_ _0492_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput7 scale[4] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_4
X_0976_ count\[24\] _0480_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0830_ true_scale\[6\] count\[5\] VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0692_ _0203_ _0214_ _0193_ _0195_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__o2bb2a_1
X_0761_ _0260_ _0278_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0959_ count\[18\] _0468_ _0447_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__o21ai_1
Xinput10 scale[7] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_4
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0813_ net16 _0344_ _0345_ _0346_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__o31ai_1
X_0675_ _0193_ _0195_ _0216_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__o21ai_1
X_0744_ true_scale\[20\] _0281_ _0067_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__mux2_1
X_1012_ net18 _0009_ VGND VGND VPWR VPWR true_scale\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0727_ _0260_ _0264_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0658_ true_scale\[15\] _0200_ _0067_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_1
X_0589_ _0120_ _0133_ _0134_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__or3_1
X_0512_ net14 true_scale\[5\] net15 VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__mux2_1
Xfanout18 net19 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0992_ count\[29\] VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 scale[5] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
X_0975_ _0482_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
X_0760_ _0294_ _0296_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__xnor2_1
X_0691_ _0154_ _0177_ _0196_ _0215_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__nor4_1
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0958_ count\[16\] count\[17\] count\[18\] _0465_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__and4_2
X_0889_ true_scale\[24\] _0061_ true_scale\[25\] VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_6_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0743_ _0278_ _0280_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__xnor2_1
X_0812_ true_scale\[24\] net16 VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__nand2_1
X_0674_ _0196_ _0199_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__or2b_1
X_1011_ net1 _0008_ VGND VGND VPWR VPWR true_scale\[13\] sky130_fd_sc_hd__dfxtp_1
X_0726_ _0260_ _0264_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__or2_1
X_0657_ _0196_ _0199_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__xnor2_1
X_0588_ _0100_ _0116_ _0115_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0511_ _0064_ VGND VGND VPWR VPWR clk_out sky130_fd_sc_hd__clkbuf_4
Xfanout19 net1 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
X_0709_ true_scale\[18\] _0248_ _0067_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_35_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0991_ _0493_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 scale[6] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_4
X_0974_ _0480_ _0481_ _0432_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__and3b_1
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0690_ _0103_ _0123_ _0133_ _0134_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_38_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0957_ _0470_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
X_0888_ _0413_ _0415_ _0416_ _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0742_ _0260_ _0264_ _0279_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a21oi_1
X_0673_ _0203_ _0214_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__xnor2_2
X_0811_ _0337_ _0334_ _0343_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1010_ net19 _0007_ VGND VGND VPWR VPWR true_scale\[12\] sky130_fd_sc_hd__dfxtp_1
X_0656_ _0155_ _0197_ _0198_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__a21oi_1
X_0725_ _0236_ _0261_ _0263_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0587_ _0122_ _0132_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0510_ net22 signal_clk_out _0063_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0639_ net6 net13 net9 VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0708_ _0245_ _0247_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0990_ _0437_ _0491_ _0492_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0973_ count\[22\] _0477_ count\[23\] VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0956_ _0468_ _0469_ _0437_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__and3b_1
XFILLER_0_27_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0887_ count\[23\] _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0810_ _0337_ _0334_ _0343_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__and3_1
X_0672_ _0204_ _0213_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__xor2_2
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0741_ _0257_ _0259_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__nor2_1
X_0939_ _0458_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0655_ _0159_ _0176_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__and2_1
X_0586_ _0129_ _0131_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__xnor2_1
X_0724_ _0240_ _0244_ _0262_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0707_ _0227_ _0229_ _0246_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__o21ai_1
X_0638_ _0145_ _0160_ _0161_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__o21bai_4
X_0569_ _0105_ _0098_ _0114_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__or3b_1
XFILLER_0_29_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0972_ count\[22\] count\[23\] _0477_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0955_ count\[16\] _0465_ count\[17\] VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__a21o_1
X_0886_ true_scale\[24\] _0061_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0740_ _0275_ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__xor2_1
X_0671_ _0211_ _0212_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__xnor2_2
X_0938_ _0456_ _0457_ _0437_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__and3b_1
X_0869_ _0398_ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0723_ _0240_ _0244_ _0227_ _0229_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__o2bb2a_1
X_0654_ _0150_ _0153_ _0159_ _0176_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__o22a_1
X_0585_ _0107_ _0113_ _0130_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0706_ _0230_ _0236_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__or2b_1
X_0637_ _0180_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__clkbuf_1
X_0568_ _0105_ _0098_ _0114_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0971_ count\[22\] _0477_ _0479_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0954_ count\[16\] count\[17\] _0465_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__and3_1
X_0885_ _0061_ _0414_ count\[22\] VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0670_ _0185_ _0188_ _0187_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_26_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0937_ count\[10\] _0453_ count\[11\] VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__a21o_1
X_0868_ true_scale\[18\] _0058_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__and2_1
X_0799_ _0322_ _0323_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0653_ _0193_ _0195_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__xnor2_2
X_0722_ _0230_ _0245_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__nor2_1
X_0584_ _0109_ _0112_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0636_ true_scale\[14\] _0179_ _0067_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_29_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0705_ _0240_ _0244_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_13_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0567_ _0107_ _0113_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0619_ net10 _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__xnor2_2
X_0970_ count\[22\] _0477_ _0433_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0953_ count\[16\] _0465_ _0467_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__a21oi_1
X_0884_ count\[22\] _0061_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0936_ count\[10\] count\[11\] _0453_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0867_ true_scale\[18\] _0058_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__nor2_1
X_0798_ _0331_ _0332_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0583_ _0123_ _0128_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__xnor2_1
X_0652_ _0139_ _0175_ _0194_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__a21oi_2
X_0721_ _0257_ _0259_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__xor2_1
X_0919_ _0443_ _0444_ _0437_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__and3b_1
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0635_ _0177_ _0178_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__xnor2_1
X_0704_ _0122_ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__xor2_2
X_0566_ _0109_ _0112_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1049_ net21 _0046_ VGND VGND VPWR VPWR count\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0618_ _0160_ _0161_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__nor2_1
X_0549_ _0095_ _0096_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0952_ count\[16\] _0465_ _0433_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__o21ai_1
X_0883_ true_scale\[23\] _0060_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0935_ count\[10\] _0453_ _0455_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a21oi_1
X_0866_ count\[16\] _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__xor2_1
X_0797_ _0330_ _0325_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0720_ _0122_ _0243_ _0258_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__o21a_1
X_0651_ _0172_ _0174_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__and2_1
X_0582_ _0126_ _0127_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0918_ count\[4\] _0355_ count\[5\] VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__a21o_1
X_0849_ _0378_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__nor2_1
X_0703_ _0241_ _0242_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0634_ _0150_ _0153_ _0155_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0565_ _0110_ _0111_ _0093_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1048_ net21 _0045_ VGND VGND VPWR VPWR count\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0617_ net7 net13 net9 VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__and3_1
X_0548_ _0079_ _0082_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__or2_2
XFILLER_0_31_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0951_ _0465_ _0466_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__nor2_1
X_0882_ _0404_ _0407_ _0409_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0934_ count\[10\] _0453_ _0433_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__o21ai_1
X_0865_ _0058_ _0395_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__nand2_1
X_0796_ _0325_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0650_ _0181_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__xnor2_2
X_0581_ net14 _0071_ _0092_ _0108_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0917_ count\[4\] count\[5\] _0355_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__and3_1
X_0848_ true_scale\[12\] _0056_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__and2_1
X_0779_ _0291_ _0306_ _0313_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__nand3_1
X_0633_ _0159_ _0176_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__xnor2_1
X_0702_ _0221_ _0107_ _0220_ _0095_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a22o_1
X_0564_ net13 _0081_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__xnor2_4
X_1047_ net20 _0044_ VGND VGND VPWR VPWR count\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0616_ net7 net13 net9 VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0547_ _0092_ _0094_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0950_ count\[15\] _0462_ _0447_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__o21ai_1
X_0881_ count\[21\] _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0795_ _0328_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0933_ _0453_ _0454_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__nor2_1
X_0864_ true_scale\[15\] true_scale\[16\] _0057_ true_scale\[17\] VGND VGND VPWR VPWR
+ _0395_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0580_ _0111_ _0125_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0916_ count\[4\] _0355_ _0442_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0847_ true_scale\[12\] _0056_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__nor2_1
X_0778_ _0291_ _0306_ _0313_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0632_ _0139_ _0175_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__xnor2_1
X_0701_ _0113_ _0123_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__xnor2_2
X_0563_ net14 _0071_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__nand2_1
X_1046_ net20 _0043_ VGND VGND VPWR VPWR count\[21\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_8_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0615_ _0139_ _0149_ _0158_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__a21boi_2
X_0546_ net14 _0071_ _0093_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1029_ net17 _0026_ VGND VGND VPWR VPWR count\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0529_ net4 net14 net5 VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ _0060_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0932_ count\[9\] _0450_ _0447_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0794_ _0204_ _0327_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0863_ _0384_ _0387_ _0391_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_21_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire11 _0232_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0915_ count\[4\] _0355_ _0433_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__o21ai_1
X_0777_ _0181_ _0312_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__xor2_1
X_0846_ count\[10\] _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__xor2_1
X_0700_ _0205_ _0226_ _0239_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__a21o_1
X_0631_ _0172_ _0174_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__xor2_1
X_0562_ _0092_ _0108_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__xnor2_4
X_1045_ net20 _0042_ VGND VGND VPWR VPWR count\[20\] sky130_fd_sc_hd__dfxtp_1
X_0829_ _0357_ _0358_ count\[6\] VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0614_ _0144_ _0148_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__nand2_1
X_0545_ net4 net5 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__nor2_1
X_1028_ net17 _0025_ VGND VGND VPWR VPWR count\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0528_ true_scale\[8\] net15 _0076_ _0077_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0931_ count\[7\] count\[8\] count\[9\] _0446_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__and4_2
X_0862_ count\[15\] _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__xnor2_1
X_0793_ _0327_ _0204_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0914_ _0441_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
X_0845_ _0056_ _0375_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__nand2_1
X_0776_ _0310_ _0311_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0630_ _0146_ _0143_ _0173_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a21bo_1
X_0561_ _0071_ _0070_ _0079_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__a21o_1
X_1044_ net20 _0041_ VGND VGND VPWR VPWR count\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0828_ count\[6\] _0357_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__and3_1
X_0759_ _0139_ _0274_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0613_ _0068_ _0155_ _0156_ _0157_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a31o_1
X_0544_ net13 _0081_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__xor2_4
X_1027_ net17 _0024_ VGND VGND VPWR VPWR count\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0527_ net6 _0075_ net15 VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0792_ _0307_ _0326_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__xor2_1
X_0930_ _0452_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
X_0861_ true_scale\[16\] _0388_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0775_ _0286_ _0289_ _0309_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__a21oi_1
X_0913_ _0355_ _0437_ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__and3b_1
X_0844_ true_scale\[9\] true_scale\[10\] _0055_ true_scale\[11\] VGND VGND VPWR VPWR
+ _0375_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0560_ net9 _0106_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__xor2_4
X_1043_ net21 _0040_ VGND VGND VPWR VPWR count\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0827_ true_scale\[5\] true_scale\[6\] true_scale\[7\] VGND VGND VPWR VPWR _0358_
+ sky130_fd_sc_hd__o21ai_1
X_0758_ _0273_ _0271_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__and2b_1
X_0689_ _0227_ _0229_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0612_ true_scale\[13\] net15 VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__and2_1
X_0543_ _0087_ _0088_ _0091_ net15 true_scale\[9\] VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a32o_1
X_1026_ net17 _0023_ VGND VGND VPWR VPWR count\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0526_ net6 _0075_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ net19 _0006_ VGND VGND VPWR VPWR true_scale\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0509_ true_scale\[26\] _0062_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0791_ net13 net10 VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__xor2_1
X_0860_ count\[14\] _0390_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ count\[28\] _0489_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0912_ count\[0\] count\[1\] count\[2\] count\[3\] VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__a31o_1
X_0774_ _0286_ _0289_ _0309_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__and3_1
X_0843_ _0363_ _0367_ _0371_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1042_ net21 _0039_ VGND VGND VPWR VPWR count\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0688_ _0204_ _0213_ _0228_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a21oi_2
X_0826_ true_scale\[5\] true_scale\[6\] true_scale\[7\] VGND VGND VPWR VPWR _0357_
+ sky130_fd_sc_hd__or3_1
X_0757_ _0139_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0611_ _0136_ _0154_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__nand2_1
X_0542_ net15 _0090_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__nor2_1
X_1025_ net17 _0022_ VGND VGND VPWR VPWR count\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_28_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0809_ _0341_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__or2_1
XANTENNA_1 _0163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0525_ _0074_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__buf_2
XFILLER_0_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1008_ net19 _0005_ VGND VGND VPWR VPWR true_scale\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0508_ true_scale\[24\] true_scale\[25\] _0061_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0790_ _0181_ _0324_ _0311_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ count\[28\] _0489_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0911_ _0439_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
X_0842_ count\[9\] _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__xnor2_1
X_0773_ _0307_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ net21 _0038_ VGND VGND VPWR VPWR count\[16\] sky130_fd_sc_hd__dfxtp_1
X_0825_ count\[4\] true_scale\[5\] _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a21bo_1
X_0756_ _0291_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__and2_1
X_0687_ _0212_ _0211_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0610_ _0136_ _0154_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__or2_1
X_0541_ _0079_ _0089_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__and2_1
X_1024_ net23 _0021_ VGND VGND VPWR VPWR true_scale\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0808_ _0338_ _0339_ _0340_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__nor3b_1
X_0739_ _0139_ _0256_ _0276_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0524_ net4 net14 net5 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_194 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1007_ net19 _0004_ VGND VGND VPWR VPWR true_scale\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0507_ true_scale\[23\] _0060_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__or2_2
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ _0489_ _0490_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0772_ net7 _0185_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__or2_1
X_0910_ _0436_ _0437_ _0438_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__and3_1
X_0841_ true_scale\[10\] _0368_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1040_ net18 _0037_ VGND VGND VPWR VPWR count\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0824_ count\[0\] count\[1\] count\[3\] count\[2\] VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__and4_2
X_0755_ _0283_ _0284_ _0290_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__or3_1
X_0686_ _0205_ _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0540_ net6 net7 VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__and2_1
X_1023_ net23 _0020_ VGND VGND VPWR VPWR true_scale\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0738_ _0255_ _0254_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__or2b_1
X_0807_ _0338_ _0339_ _0340_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0669_ _0207_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__xor2_2
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0523_ _0073_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__clkbuf_1
X_1006_ net19 _0003_ VGND VGND VPWR VPWR true_scale\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0506_ true_scale\[21\] true_scale\[22\] _0059_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ count\[27\] _0486_ _0447_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0771_ net7 _0185_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__nand2_1
X_0840_ count\[8\] _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ _0477_ _0478_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0823_ _0354_ _0352_ _0068_ true_scale\[26\] VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__o2bb2a_1
X_0685_ _0223_ _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__xor2_2
X_0754_ _0283_ _0284_ _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1022_ net22 _0019_ VGND VGND VPWR VPWR true_scale\[24\] sky130_fd_sc_hd__dfxtp_1
X_0806_ net7 _0185_ _0326_ _0328_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__a31o_1
X_0737_ _0139_ _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__xnor2_2
X_0668_ _0096_ _0209_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0599_ _0123_ _0143_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0522_ true_scale\[7\] _0072_ _0068_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_16_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1005_ net19 _0002_ VGND VGND VPWR VPWR true_scale\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0505_ true_scale\[18\] true_scale\[19\] true_scale\[20\] _0058_ VGND VGND VPWR VPWR
+ _0059_ sky130_fd_sc_hd__or4_2
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_26U9NK c1_n3146_n1500# m3_n3186_n1540#
X0 c1_n3146_n1500# m3_n3186_n1540# sky130_fd_pr__cap_mim_m3_1 l=15 w=30
.ends

.subckt sky130_fd_pr__pfet_01v8_AXJJQ9 a_158_n197# a_n874_n197# a_n416_n100# a_874_n100#
+ w_n968_n200# a_n358_n197# a_358_n100# a_416_n197# a_n100_n197# a_100_n100# a_n674_n100#
+ a_n158_n100# a_n616_n197# a_674_n197# a_616_n100# a_n932_n100#
X0 a_874_n100# a_674_n197# a_616_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1 a_n158_n100# a_n358_n197# a_n416_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 a_100_n100# a_n100_n197# a_n158_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3 a_n674_n100# a_n874_n197# a_n932_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X4 a_616_n100# a_416_n197# a_358_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X5 a_358_n100# a_158_n197# a_100_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X6 a_n416_n100# a_n616_n197# a_n674_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_HD5U9F a_n129_n150# a_n221_n150# a_63_n150# a_111_172#
+ a_n33_n150# a_n81_172# a_159_n150# a_15_n238# a_n177_n238# VSUBS
X0 a_159_n150# a_111_172# a_63_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.465 pd=3.62 as=0.248 ps=1.83 w=1.5 l=0.15
X1 a_63_n150# a_15_n238# a_n33_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.248 ps=1.83 w=1.5 l=0.15
X2 a_n129_n150# a_n177_n238# a_n221_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.465 ps=3.62 w=1.5 l=0.15
X3 a_n33_n150# a_n81_172# a_n129_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.248 pd=1.83 as=0.248 ps=1.83 w=1.5 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_5VPKLS a_n29_n100# a_487_n100# a_n229_n188# a_287_n188#
+ a_n287_n100# a_n487_n188# a_229_n100# a_n545_n100# a_29_n188# VSUBS
X0 a_n287_n100# a_n487_n188# a_n545_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1 a_n29_n100# a_n229_n188# a_n287_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 a_229_n100# a_29_n188# a_n29_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3 a_487_n100# a_287_n188# a_229_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_99C25S a_n229_n1597# a_n545_n1500# a_n29_n1500# a_229_n1500#
+ a_287_n1597# a_29_n1597# a_n487_n1597# a_487_n1500# a_n287_n1500# w_n581_n1600#
X0 a_487_n1500# a_287_n1597# a_229_n1500# w_n581_n1600# sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.6 as=2.17 ps=15.3 w=15 l=1
X1 a_n287_n1500# a_n487_n1597# a_n545_n1500# w_n581_n1600# sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=4.35 ps=30.6 w=15 l=1
X2 a_n29_n1500# a_n229_n1597# a_n287_n1500# w_n581_n1600# sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
X3 a_229_n1500# a_29_n1597# a_n29_n1500# w_n581_n1600# sky130_fd_pr__pfet_01v8 ad=2.17 pd=15.3 as=2.17 ps=15.3 w=15 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_MMM6UU a_n287_n500# a_n487_n588# a_745_n500# a_545_n588#
+ a_229_n500# a_n545_n500# a_29_n588# a_n745_n588# a_n29_n500# a_487_n500# a_n229_n588#
+ a_287_n588# a_n803_n500# VSUBS
X0 a_487_n500# a_287_n588# a_229_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_745_n500# a_545_n588# a_487_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=1
X2 a_n29_n500# a_n229_n588# a_n287_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_229_n500# a_29_n588# a_n29_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_n545_n500# a_n745_n588# a_n803_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=1
X5 a_n287_n500# a_n487_n588# a_n545_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt buffer vd ib out in gnd
Xsky130_fd_pr__cap_mim_m3_1_26U9NK_0 out d sky130_fd_pr__cap_mim_m3_1_26U9NK
Xsky130_fd_pr__pfet_01v8_AXJJQ9_0 a vd a a vd a vd a a a vd vd a a a vd sky130_fd_pr__pfet_01v8_AXJJQ9
Xsky130_fd_pr__pfet_01v8_AXJJQ9_1 b b vd vd vd b b b b vd b b b vd vd b sky130_fd_pr__pfet_01v8_AXJJQ9
Xsky130_fd_pr__nfet_01v8_HD5U9F_1 a a b b c out b in a gnd sky130_fd_pr__nfet_01v8_HD5U9F
Xsky130_fd_pr__nfet_01v8_5VPKLS_0 gnd c ib c ib ib c ib ib gnd sky130_fd_pr__nfet_01v8_5VPKLS
Xsky130_fd_pr__pfet_01v8_99C25S_0 a d vd d d a d d d vd sky130_fd_pr__pfet_01v8_99C25S
Xsky130_fd_pr__pfet_01v8_99C25S_1 b out vd out out b out out out vd sky130_fd_pr__pfet_01v8_99C25S
XXM10 d d gnd gnd out gnd d gnd gnd gnd d d gnd gnd sky130_fd_pr__nfet_01v8_MMM6UU
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_XMXTTL a_546_450# a_n118_450# a_546_n882#
+ a_n450_450# a_n450_n882# a_n284_n882# a_n118_n882# a_n616_450# a_380_n882# a_48_450#
+ a_380_450# a_n616_n882# a_214_n882# a_214_450# a_n284_450# a_48_n882# VSUBS
X0 a_n616_450# a_n616_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X1 a_380_450# a_380_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X2 a_546_450# a_546_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X3 a_214_450# a_214_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X4 a_n284_450# a_n284_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X5 a_n450_450# a_n450_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X6 a_48_450# a_48_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.5
X7 a_n118_450# a_n118_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.5
.ends

.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.213 ps=1.67 w=1 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3 VPWR a_1283_21# a_1847_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9 Q_N a_1847_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_1283_21# a_1847_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X12 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X13 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X17 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X18 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X19 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X20 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X26 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X27 Q_N a_1847_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X28 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X29 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X31 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_XGSNAL a_n33_n397# a_n73_n300# a_15_n300# w_n211_n519#
X0 a_15_n300# a_n33_n397# a_n73_n300# w_n211_n519# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_QABHPF a_546_200# a_n118_200# a_546_n632#
+ a_n450_200# a_n450_n632# a_n284_n632# a_n118_n632# a_n616_200# a_48_200# a_380_n632#
+ a_380_200# a_n616_n632# a_214_n632# a_214_200# a_n284_200# a_48_n632# VSUBS
X0 a_n450_200# a_n450_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2
X1 a_n118_200# a_n118_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2
X2 a_n616_200# a_n616_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2
X3 a_380_200# a_380_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2
X4 a_546_200# a_546_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2
X5 a_214_200# a_214_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2
X6 a_n284_200# a_n284_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2
X7 a_48_200# a_48_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_A4KLY5 c1_n2866_n2720# m3_n2906_n2760#
X0 c1_n2866_n2720# m3_n2906_n2760# sky130_fd_pr__cap_mim_m3_1 l=27.2 w=27.2
.ends

.subckt sigma-delta out vpwr clk reset_b_dff gnd vd in
Xsky130_fd_pr__res_xhigh_po_0p35_XMXTTL_1 m1_n1920_4820# m1_n2580_4820# in_int m1_n2940_4820#
+ m1_n2760_3480# m1_n2760_3480# m1_n2420_3480# m1_n2940_4820# m1_n2100_3480# m1_n2260_4820#
+ m1_n1920_4820# in m1_n2100_3480# m1_n2260_4820# m1_n2580_4820# m1_n2420_3480# gnd
+ sky130_fd_pr__res_xhigh_po_0p35_XMXTTL
Xx1 clk x1/D reset_b_dff gnd gnd vpwr vpwr x1/Q out sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_pr__res_xhigh_po_0p35_XMXTTL_2 m1_n440_4820# m1_n1100_4820# x1/Q m1_n1440_4820#
+ m1_n1260_3480# m1_n1260_3480# m1_n940_3480# m1_n1440_4820# m1_n620_3480# m1_n780_4820#
+ m1_n440_4820# in_int m1_n620_3480# m1_n780_4820# m1_n1100_4820# m1_n940_3480# gnd
+ sky130_fd_pr__res_xhigh_po_0p35_XMXTTL
Xsky130_fd_pr__nfet_01v8_648S5X_0 x1/D in_comp gnd gnd sky130_fd_pr__nfet_01v8_648S5X
XXP1 in_comp x1/D vd vd sky130_fd_pr__pfet_01v8_XGSNAL
Xsky130_fd_pr__res_xhigh_po_0p35_QABHPF_0 in_comp m1_n2360_2660# m1_n1860_1820# m1_n2700_2660#
+ m1_n2860_1820# m1_n2520_1820# m1_n2520_1820# in_int m1_n2360_2660# m1_n1860_1820#
+ m1_n2040_2660# m1_n2860_1820# m1_n2200_1820# m1_n2040_2660# m1_n2700_2660# m1_n2200_1820#
+ gnd sky130_fd_pr__res_xhigh_po_0p35_QABHPF
Xsky130_fd_pr__cap_mim_m3_1_A4KLY5_0 in_comp gnd sky130_fd_pr__cap_mim_m3_1_A4KLY5
Xsky130_fd_pr__cap_mim_m3_1_A4KLY5_1 in_int gnd sky130_fd_pr__cap_mim_m3_1_A4KLY5
.ends

.subckt tt_um_hugodiasg_temp-sensor_clock-divider clk ena rst_n ua[0] ua[1] ua[2]
+ ua[3] ua[4] ua[5] ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5]
+ ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6]
+ uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6]
+ uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6]
+ uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] VDPWR VGND
Xsensor_0 VDPWR ua[4] ua[5] VGND sensor
Xclock_divider_0 clk uo_out[0] rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4]
+ ui_in[5] ui_in[6] ui_in[7] VDPWR VGND clock_divider
Xbuffer_0 VDPWR ua[2] ua[1] ua[3] VGND buffer
Xsigma-delta_0 uo_out[7] VDPWR clk VDPWR VGND VDPWR ua[0] sigma-delta
.ends

