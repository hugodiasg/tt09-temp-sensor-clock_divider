MACRO clock_divider
  CLASS BLOCK ;
  FOREIGN clock_divider ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.580 2.480 23.180 117.200 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 117.200 ;
    END
  END VPWR
  PIN clk_in
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 118.000 19.080 120.000 19.680 ;
    END
  END clk_in
  PIN clk_out
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 118.000 97.960 120.000 98.560 ;
    END
  END clk_out
  PIN nrst
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 118.000 58.520 120.000 59.120 ;
    END
  END nrst
  PIN scale[0]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 8.370 118.000 8.650 120.000 ;
    END
  END scale[0]
  PIN scale[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 23.090 118.000 23.370 120.000 ;
    END
  END scale[1]
  PIN scale[2]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 37.810 118.000 38.090 120.000 ;
    END
  END scale[2]
  PIN scale[3]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 52.530 118.000 52.810 120.000 ;
    END
  END scale[3]
  PIN scale[4]
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 67.250 118.000 67.530 120.000 ;
    END
  END scale[4]
  PIN scale[5]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.970 118.000 82.250 120.000 ;
    END
  END scale[5]
  PIN scale[6]
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 118.000 96.970 120.000 ;
    END
  END scale[6]
  PIN scale[7]
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 111.410 118.000 111.690 120.000 ;
    END
  END scale[7]
  OBS
      LAYER nwell ;
        RECT 2.570 2.635 117.030 117.045 ;
      LAYER li1 ;
        RECT 2.760 2.635 116.840 117.045 ;
      LAYER met1 ;
        RECT 2.760 2.480 116.840 117.200 ;
      LAYER met2 ;
        RECT 8.930 117.720 22.810 118.730 ;
        RECT 23.650 117.720 37.530 118.730 ;
        RECT 38.370 117.720 52.250 118.730 ;
        RECT 53.090 117.720 66.970 118.730 ;
        RECT 67.810 117.720 81.690 118.730 ;
        RECT 82.530 117.720 96.410 118.730 ;
        RECT 97.250 117.720 111.130 118.730 ;
        RECT 111.970 117.720 115.370 118.730 ;
        RECT 8.380 2.535 115.370 117.720 ;
      LAYER met3 ;
        RECT 18.290 98.960 118.000 117.125 ;
        RECT 18.290 97.560 117.600 98.960 ;
        RECT 18.290 59.520 118.000 97.560 ;
        RECT 18.290 58.120 117.600 59.520 ;
        RECT 18.290 20.080 118.000 58.120 ;
        RECT 18.290 18.680 117.600 20.080 ;
        RECT 18.290 2.555 118.000 18.680 ;
  END
END clock_divider
END LIBRARY

