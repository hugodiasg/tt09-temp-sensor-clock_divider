magic
tech sky130A
magscale 1 2
timestamp 1729285596
<< viali >>
rect 1961 23273 1995 23307
rect 7849 23273 7883 23307
rect 19257 23273 19291 23307
rect 10425 23205 10459 23239
rect 13829 23205 13863 23239
rect 19533 23205 19567 23239
rect 19901 23205 19935 23239
rect 21557 23205 21591 23239
rect 1777 23137 1811 23171
rect 4721 23137 4755 23171
rect 6101 23137 6135 23171
rect 6285 23137 6319 23171
rect 7573 23137 7607 23171
rect 7757 23137 7791 23171
rect 8033 23137 8067 23171
rect 11069 23137 11103 23171
rect 11161 23137 11195 23171
rect 11345 23137 11379 23171
rect 11437 23137 11471 23171
rect 13553 23137 13587 23171
rect 16497 23137 16531 23171
rect 18981 23137 19015 23171
rect 19993 23137 20027 23171
rect 20177 23137 20211 23171
rect 21281 23137 21315 23171
rect 21373 23137 21407 23171
rect 21649 23137 21683 23171
rect 21741 23137 21775 23171
rect 21925 23137 21959 23171
rect 22385 23137 22419 23171
rect 18797 23069 18831 23103
rect 19349 23069 19383 23103
rect 22569 23069 22603 23103
rect 5917 23001 5951 23035
rect 10609 23001 10643 23035
rect 4905 22933 4939 22967
rect 6469 22933 6503 22967
rect 7665 22933 7699 22967
rect 11621 22933 11655 22967
rect 16681 22933 16715 22967
rect 19993 22933 20027 22967
rect 21465 22933 21499 22967
rect 21925 22933 21959 22967
rect 5089 22729 5123 22763
rect 9873 22729 9907 22763
rect 13185 22729 13219 22763
rect 14289 22729 14323 22763
rect 15301 22729 15335 22763
rect 18337 22729 18371 22763
rect 18521 22729 18555 22763
rect 20729 22729 20763 22763
rect 21557 22729 21591 22763
rect 5549 22661 5583 22695
rect 10149 22661 10183 22695
rect 12817 22661 12851 22695
rect 14105 22661 14139 22695
rect 15485 22661 15519 22695
rect 16497 22661 16531 22695
rect 21833 22661 21867 22695
rect 9413 22593 9447 22627
rect 11345 22593 11379 22627
rect 11529 22593 11563 22627
rect 13093 22593 13127 22627
rect 13553 22593 13587 22627
rect 13737 22593 13771 22627
rect 15853 22593 15887 22627
rect 19257 22593 19291 22627
rect 19993 22593 20027 22627
rect 21097 22593 21131 22627
rect 5365 22525 5399 22559
rect 5457 22525 5491 22559
rect 5733 22525 5767 22559
rect 6377 22525 6411 22559
rect 7205 22525 7239 22559
rect 8401 22525 8435 22559
rect 9229 22525 9263 22559
rect 10425 22525 10459 22559
rect 11253 22525 11287 22559
rect 11621 22525 11655 22559
rect 11713 22525 11747 22559
rect 11897 22525 11931 22559
rect 11989 22525 12023 22559
rect 12173 22525 12207 22559
rect 12541 22525 12575 22559
rect 12633 22525 12667 22559
rect 13277 22525 13311 22559
rect 13369 22525 13403 22559
rect 14013 22525 14047 22559
rect 14565 22525 14599 22559
rect 14658 22525 14692 22559
rect 15945 22525 15979 22559
rect 16221 22525 16255 22559
rect 19809 22525 19843 22559
rect 21189 22525 21223 22559
rect 14243 22491 14277 22525
rect 18383 22491 18417 22525
rect 4905 22457 4939 22491
rect 6193 22457 6227 22491
rect 9689 22457 9723 22491
rect 10149 22457 10183 22491
rect 10333 22457 10367 22491
rect 12817 22457 12851 22491
rect 14473 22457 14507 22491
rect 15117 22457 15151 22491
rect 16497 22457 16531 22491
rect 16773 22457 16807 22491
rect 17509 22457 17543 22491
rect 17601 22457 17635 22491
rect 17785 22457 17819 22491
rect 18153 22457 18187 22491
rect 18705 22457 18739 22491
rect 18889 22457 18923 22491
rect 20545 22457 20579 22491
rect 20761 22457 20795 22491
rect 22109 22457 22143 22491
rect 5089 22389 5123 22423
rect 8493 22389 8527 22423
rect 9045 22389 9079 22423
rect 9889 22389 9923 22423
rect 10057 22389 10091 22423
rect 10885 22389 10919 22423
rect 13921 22389 13955 22423
rect 14933 22389 14967 22423
rect 15317 22389 15351 22423
rect 15577 22389 15611 22423
rect 16313 22389 16347 22423
rect 17969 22389 18003 22423
rect 19073 22389 19107 22423
rect 20913 22389 20947 22423
rect 21649 22389 21683 22423
rect 12725 22185 12759 22219
rect 15485 22185 15519 22219
rect 18337 22185 18371 22219
rect 18629 22185 18663 22219
rect 18797 22185 18831 22219
rect 10701 22117 10735 22151
rect 15577 22117 15611 22151
rect 15945 22117 15979 22151
rect 18429 22117 18463 22151
rect 21281 22117 21315 22151
rect 22569 22117 22603 22151
rect 5457 22049 5491 22083
rect 5917 22049 5951 22083
rect 6285 22049 6319 22083
rect 6561 22049 6595 22083
rect 7757 22049 7791 22083
rect 8493 22049 8527 22083
rect 8861 22049 8895 22083
rect 9045 22049 9079 22083
rect 9597 22049 9631 22083
rect 10333 22049 10367 22083
rect 10517 22049 10551 22083
rect 11161 22049 11195 22083
rect 11437 22049 11471 22083
rect 11805 22049 11839 22083
rect 12081 22049 12115 22083
rect 12265 22049 12299 22083
rect 12357 22049 12391 22083
rect 12449 22049 12483 22083
rect 13185 22049 13219 22083
rect 14105 22049 14139 22083
rect 15761 22049 15795 22083
rect 16129 22049 16163 22083
rect 16589 22049 16623 22083
rect 16957 22049 16991 22083
rect 17417 22049 17451 22083
rect 17509 22049 17543 22083
rect 17686 22049 17720 22083
rect 17969 22049 18003 22083
rect 19073 22049 19107 22083
rect 19717 22049 19751 22083
rect 19993 22049 20027 22083
rect 20913 22049 20947 22083
rect 21373 22049 21407 22083
rect 21557 22049 21591 22083
rect 21649 22049 21683 22083
rect 21925 22049 21959 22083
rect 22293 22049 22327 22083
rect 22385 22049 22419 22083
rect 9321 21981 9355 22015
rect 10241 21981 10275 22015
rect 11989 21981 12023 22015
rect 13093 21981 13127 22015
rect 13829 21981 13863 22015
rect 14749 21981 14783 22015
rect 15025 21981 15059 22015
rect 15117 21981 15151 22015
rect 17601 21981 17635 22015
rect 18061 21981 18095 22015
rect 22017 21981 22051 22015
rect 22753 21981 22787 22015
rect 6009 21913 6043 21947
rect 7481 21913 7515 21947
rect 8953 21913 8987 21947
rect 5273 21845 5307 21879
rect 11897 21845 11931 21879
rect 12909 21845 12943 21879
rect 14841 21845 14875 21879
rect 18613 21845 18647 21879
rect 19257 21845 19291 21879
rect 20545 21845 20579 21879
rect 21741 21845 21775 21879
rect 22109 21845 22143 21879
rect 22201 21845 22235 21879
rect 16773 21641 16807 21675
rect 21465 21641 21499 21675
rect 5273 21573 5307 21607
rect 6285 21573 6319 21607
rect 8125 21573 8159 21607
rect 9597 21573 9631 21607
rect 10241 21573 10275 21607
rect 10885 21573 10919 21607
rect 13369 21573 13403 21607
rect 15577 21573 15611 21607
rect 17325 21573 17359 21607
rect 18245 21573 18279 21607
rect 19625 21573 19659 21607
rect 21833 21573 21867 21607
rect 22109 21573 22143 21607
rect 6009 21505 6043 21539
rect 7205 21505 7239 21539
rect 7665 21505 7699 21539
rect 8861 21505 8895 21539
rect 9045 21505 9079 21539
rect 9229 21505 9263 21539
rect 9689 21505 9723 21539
rect 12081 21505 12115 21539
rect 14657 21505 14691 21539
rect 16037 21505 16071 21539
rect 16589 21505 16623 21539
rect 18981 21505 19015 21539
rect 19257 21505 19291 21539
rect 22017 21505 22051 21539
rect 5917 21437 5951 21471
rect 7757 21437 7791 21471
rect 9781 21437 9815 21471
rect 10057 21437 10091 21471
rect 10425 21437 10459 21471
rect 10701 21437 10735 21471
rect 11069 21437 11103 21471
rect 12448 21437 12482 21471
rect 12541 21437 12575 21471
rect 13093 21437 13127 21471
rect 13185 21437 13219 21471
rect 13369 21437 13403 21471
rect 13921 21437 13955 21471
rect 14013 21437 14047 21471
rect 14749 21437 14783 21471
rect 15945 21437 15979 21471
rect 16497 21437 16531 21471
rect 17141 21437 17175 21471
rect 17693 21437 17727 21471
rect 17877 21437 17911 21471
rect 17969 21437 18003 21471
rect 18061 21437 18095 21471
rect 18245 21437 18279 21471
rect 18521 21437 18555 21471
rect 18889 21437 18923 21471
rect 19349 21437 19383 21471
rect 20575 21437 20609 21471
rect 20729 21437 20763 21471
rect 21005 21437 21039 21471
rect 21097 21437 21131 21471
rect 21281 21437 21315 21471
rect 22109 21437 22143 21471
rect 22293 21437 22327 21471
rect 4997 21369 5031 21403
rect 6377 21369 6411 21403
rect 8769 21369 8803 21403
rect 16957 21369 16991 21403
rect 18429 21369 18463 21403
rect 19625 21369 19659 21403
rect 21557 21369 21591 21403
rect 5457 21301 5491 21335
rect 8401 21301 8435 21335
rect 9873 21301 9907 21335
rect 10517 21301 10551 21335
rect 12173 21301 12207 21335
rect 13553 21301 13587 21335
rect 14197 21301 14231 21335
rect 15393 21301 15427 21335
rect 17509 21301 17543 21335
rect 19441 21301 19475 21335
rect 20361 21301 20395 21335
rect 10701 21097 10735 21131
rect 11253 21097 11287 21131
rect 14105 21097 14139 21131
rect 16497 21097 16531 21131
rect 17325 21097 17359 21131
rect 6469 21029 6503 21063
rect 10241 21029 10275 21063
rect 14749 21029 14783 21063
rect 4537 20961 4571 20995
rect 4997 20961 5031 20995
rect 5917 20961 5951 20995
rect 6193 20961 6227 20995
rect 6653 20961 6687 20995
rect 8217 20961 8251 20995
rect 8861 20961 8895 20995
rect 9505 20961 9539 20995
rect 9689 20961 9723 20995
rect 9781 20961 9815 20995
rect 10149 20961 10183 20995
rect 10333 20961 10367 20995
rect 10609 20961 10643 20995
rect 10793 20961 10827 20995
rect 11069 20961 11103 20995
rect 11437 20961 11471 20995
rect 13737 20961 13771 20995
rect 13921 20961 13955 20995
rect 15485 20961 15519 20995
rect 16313 20961 16347 20995
rect 16497 20961 16531 20995
rect 17233 20961 17267 20995
rect 17417 20961 17451 20995
rect 20269 20961 20303 20995
rect 20453 20961 20487 20995
rect 20545 20961 20579 20995
rect 20699 20961 20733 20995
rect 20913 20961 20947 20995
rect 21649 20961 21683 20995
rect 21741 20961 21775 20995
rect 22385 20961 22419 20995
rect 4629 20893 4663 20927
rect 4721 20893 4755 20927
rect 6101 20893 6135 20927
rect 21465 20893 21499 20927
rect 21557 20893 21591 20927
rect 5365 20825 5399 20859
rect 6009 20825 6043 20859
rect 6377 20825 6411 20859
rect 22109 20825 22143 20859
rect 4905 20757 4939 20791
rect 5457 20757 5491 20791
rect 6837 20757 6871 20791
rect 9321 20757 9355 20791
rect 11437 20757 11471 20791
rect 13737 20757 13771 20791
rect 20361 20757 20395 20791
rect 21281 20757 21315 20791
rect 21925 20757 21959 20791
rect 5089 20553 5123 20587
rect 6009 20553 6043 20587
rect 10333 20553 10367 20587
rect 14657 20553 14691 20587
rect 21281 20553 21315 20587
rect 7021 20485 7055 20519
rect 21005 20485 21039 20519
rect 5181 20417 5215 20451
rect 5641 20417 5675 20451
rect 5917 20417 5951 20451
rect 6101 20417 6135 20451
rect 13553 20417 13587 20451
rect 14289 20417 14323 20451
rect 17233 20417 17267 20451
rect 5273 20349 5307 20383
rect 5549 20349 5583 20383
rect 6009 20349 6043 20383
rect 6653 20349 6687 20383
rect 6837 20349 6871 20383
rect 6929 20349 6963 20383
rect 7113 20349 7147 20383
rect 8401 20349 8435 20383
rect 8493 20349 8527 20383
rect 8677 20349 8711 20383
rect 10333 20349 10367 20383
rect 10517 20349 10551 20383
rect 12633 20349 12667 20383
rect 12817 20349 12851 20383
rect 13737 20349 13771 20383
rect 14473 20349 14507 20383
rect 17325 20349 17359 20383
rect 17601 20349 17635 20383
rect 17694 20349 17728 20383
rect 18705 20349 18739 20383
rect 18889 20349 18923 20383
rect 20637 20349 20671 20383
rect 20729 20349 20763 20383
rect 21005 20349 21039 20383
rect 22201 20349 22235 20383
rect 20821 20281 20855 20315
rect 21097 20281 21131 20315
rect 21297 20281 21331 20315
rect 21741 20281 21775 20315
rect 4905 20213 4939 20247
rect 6377 20213 6411 20247
rect 6837 20213 6871 20247
rect 8861 20213 8895 20247
rect 13001 20213 13035 20247
rect 13921 20213 13955 20247
rect 16957 20213 16991 20247
rect 17969 20213 18003 20247
rect 18797 20213 18831 20247
rect 20453 20213 20487 20247
rect 21465 20213 21499 20247
rect 21833 20213 21867 20247
rect 22385 20213 22419 20247
rect 7389 20009 7423 20043
rect 11713 20009 11747 20043
rect 13553 20009 13587 20043
rect 18153 20009 18187 20043
rect 19241 20009 19275 20043
rect 20177 20009 20211 20043
rect 21281 20009 21315 20043
rect 6009 19941 6043 19975
rect 8861 19941 8895 19975
rect 13645 19941 13679 19975
rect 17049 19941 17083 19975
rect 19441 19941 19475 19975
rect 21925 19941 21959 19975
rect 22201 19941 22235 19975
rect 5917 19873 5951 19907
rect 6193 19873 6227 19907
rect 6653 19873 6687 19907
rect 7573 19873 7607 19907
rect 7849 19873 7883 19907
rect 8401 19873 8435 19907
rect 10333 19873 10367 19907
rect 10701 19873 10735 19907
rect 11345 19873 11379 19907
rect 12449 19873 12483 19907
rect 13185 19873 13219 19907
rect 13829 19873 13863 19907
rect 13921 19873 13955 19907
rect 14197 19873 14231 19907
rect 16957 19873 16991 19907
rect 17141 19873 17175 19907
rect 17417 19873 17451 19907
rect 18061 19873 18095 19907
rect 18337 19873 18371 19907
rect 18521 19873 18555 19907
rect 18613 19873 18647 19907
rect 19717 19873 19751 19907
rect 19809 19873 19843 19907
rect 19993 19873 20027 19907
rect 20269 19873 20303 19907
rect 20361 19873 20395 19907
rect 20545 19873 20579 19907
rect 20637 19873 20671 19907
rect 20729 19873 20763 19907
rect 20913 19873 20947 19907
rect 21097 19873 21131 19907
rect 22017 19873 22051 19907
rect 22293 19873 22327 19907
rect 22385 19873 22419 19907
rect 22661 19873 22695 19907
rect 6561 19805 6595 19839
rect 8309 19805 8343 19839
rect 11253 19805 11287 19839
rect 12357 19805 12391 19839
rect 12817 19805 12851 19839
rect 13277 19805 13311 19839
rect 14289 19805 14323 19839
rect 17325 19805 17359 19839
rect 18705 19805 18739 19839
rect 18797 19805 18831 19839
rect 18981 19805 19015 19839
rect 21649 19805 21683 19839
rect 21741 19805 21775 19839
rect 22753 19805 22787 19839
rect 6193 19737 6227 19771
rect 7021 19737 7055 19771
rect 7757 19737 7791 19771
rect 8769 19737 8803 19771
rect 13921 19737 13955 19771
rect 17785 19737 17819 19771
rect 18337 19737 18371 19771
rect 14565 19669 14599 19703
rect 19073 19669 19107 19703
rect 19257 19669 19291 19703
rect 20269 19669 20303 19703
rect 22569 19669 22603 19703
rect 22661 19669 22695 19703
rect 23029 19669 23063 19703
rect 5641 19465 5675 19499
rect 7205 19465 7239 19499
rect 8125 19465 8159 19499
rect 18521 19465 18555 19499
rect 20729 19465 20763 19499
rect 9597 19397 9631 19431
rect 16589 19397 16623 19431
rect 7757 19329 7791 19363
rect 13553 19329 13587 19363
rect 15485 19329 15519 19363
rect 15761 19329 15795 19363
rect 20177 19329 20211 19363
rect 20361 19329 20395 19363
rect 6837 19261 6871 19295
rect 7021 19261 7055 19295
rect 7849 19261 7883 19295
rect 8677 19261 8711 19295
rect 8861 19261 8895 19295
rect 9781 19261 9815 19295
rect 10425 19261 10459 19295
rect 11989 19261 12023 19295
rect 12817 19261 12851 19295
rect 13645 19261 13679 19295
rect 13829 19261 13863 19295
rect 14105 19261 14139 19295
rect 14259 19261 14293 19295
rect 14565 19261 14599 19295
rect 14749 19261 14783 19295
rect 15393 19261 15427 19295
rect 15853 19261 15887 19295
rect 16037 19261 16071 19295
rect 16313 19261 16347 19295
rect 16405 19261 16439 19295
rect 17969 19261 18003 19295
rect 18061 19261 18095 19295
rect 18337 19261 18371 19295
rect 18521 19261 18555 19295
rect 18705 19261 18739 19295
rect 18889 19261 18923 19295
rect 20269 19261 20303 19295
rect 20453 19261 20487 19295
rect 20637 19261 20671 19295
rect 21100 19261 21134 19295
rect 22486 19261 22520 19295
rect 22753 19261 22787 19295
rect 5457 19193 5491 19227
rect 14013 19193 14047 19227
rect 16221 19193 16255 19227
rect 16589 19193 16623 19227
rect 5657 19125 5691 19159
rect 5825 19125 5859 19159
rect 8861 19125 8895 19159
rect 14473 19125 14507 19159
rect 14657 19125 14691 19159
rect 18245 19125 18279 19159
rect 18797 19125 18831 19159
rect 19993 19125 20027 19159
rect 21097 19125 21131 19159
rect 21281 19125 21315 19159
rect 21373 19125 21407 19159
rect 7021 18921 7055 18955
rect 8309 18921 8343 18955
rect 9137 18921 9171 18955
rect 14289 18921 14323 18955
rect 22661 18921 22695 18955
rect 6469 18853 6503 18887
rect 10057 18853 10091 18887
rect 12081 18853 12115 18887
rect 13921 18853 13955 18887
rect 19800 18853 19834 18887
rect 21526 18853 21560 18887
rect 5273 18785 5307 18819
rect 5825 18785 5859 18819
rect 6009 18785 6043 18819
rect 6285 18785 6319 18819
rect 6837 18785 6871 18819
rect 7113 18785 7147 18819
rect 7297 18785 7331 18819
rect 7481 18785 7515 18819
rect 8861 18785 8895 18819
rect 8953 18785 8987 18819
rect 9597 18785 9631 18819
rect 9873 18785 9907 18819
rect 10609 18785 10643 18819
rect 10977 18785 11011 18819
rect 11345 18785 11379 18819
rect 11805 18785 11839 18819
rect 12357 18785 12391 18819
rect 13645 18785 13679 18819
rect 13737 18785 13771 18819
rect 14197 18785 14231 18819
rect 14473 18785 14507 18819
rect 14749 18785 14783 18819
rect 15209 18785 15243 18819
rect 15485 18785 15519 18819
rect 16497 18785 16531 18819
rect 18705 18785 18739 18819
rect 18797 18785 18831 18819
rect 18981 18785 19015 18819
rect 22845 18785 22879 18819
rect 22937 18785 22971 18819
rect 5365 18717 5399 18751
rect 6653 18717 6687 18751
rect 8493 18717 8527 18751
rect 9505 18717 9539 18751
rect 10425 18717 10459 18751
rect 12265 18717 12299 18751
rect 13921 18717 13955 18751
rect 14657 18717 14691 18751
rect 16405 18717 16439 18751
rect 18429 18717 18463 18751
rect 19533 18717 19567 18751
rect 21281 18717 21315 18751
rect 12725 18649 12759 18683
rect 14473 18649 14507 18683
rect 15669 18649 15703 18683
rect 16129 18649 16163 18683
rect 5549 18581 5583 18615
rect 9321 18581 9355 18615
rect 10241 18581 10275 18615
rect 10793 18581 10827 18615
rect 15025 18581 15059 18615
rect 15301 18581 15335 18615
rect 18521 18581 18555 18615
rect 18613 18581 18647 18615
rect 18797 18581 18831 18615
rect 20913 18581 20947 18615
rect 4445 18377 4479 18411
rect 7941 18377 7975 18411
rect 8769 18377 8803 18411
rect 10333 18377 10367 18411
rect 11621 18377 11655 18411
rect 15209 18377 15243 18411
rect 18521 18377 18555 18411
rect 20361 18377 20395 18411
rect 21097 18377 21131 18411
rect 9505 18309 9539 18343
rect 12173 18309 12207 18343
rect 19073 18309 19107 18343
rect 21557 18309 21591 18343
rect 5273 18241 5307 18275
rect 6745 18241 6779 18275
rect 7205 18241 7239 18275
rect 7297 18241 7331 18275
rect 7849 18241 7883 18275
rect 10885 18241 10919 18275
rect 11345 18241 11379 18275
rect 11805 18241 11839 18275
rect 14841 18241 14875 18275
rect 15117 18241 15151 18275
rect 16221 18241 16255 18275
rect 18981 18241 19015 18275
rect 20729 18241 20763 18275
rect 4537 18173 4571 18207
rect 5181 18173 5215 18207
rect 5917 18173 5951 18207
rect 6193 18173 6227 18207
rect 6837 18173 6871 18207
rect 7665 18173 7699 18207
rect 7941 18173 7975 18207
rect 8125 18173 8159 18207
rect 8401 18173 8435 18207
rect 8585 18173 8619 18207
rect 8953 18173 8987 18207
rect 9137 18173 9171 18207
rect 9229 18173 9263 18207
rect 9321 18173 9355 18207
rect 9597 18173 9631 18207
rect 9781 18173 9815 18207
rect 10241 18173 10275 18207
rect 10977 18173 11011 18207
rect 11621 18173 11655 18207
rect 11989 18173 12023 18207
rect 12081 18173 12115 18207
rect 12357 18173 12391 18207
rect 14749 18173 14783 18207
rect 15209 18173 15243 18207
rect 15393 18173 15427 18207
rect 16313 18173 16347 18207
rect 16773 18173 16807 18207
rect 16957 18173 16991 18207
rect 17509 18173 17543 18207
rect 17693 18173 17727 18207
rect 17877 18173 17911 18207
rect 18153 18173 18187 18207
rect 18521 18173 18555 18207
rect 18889 18173 18923 18207
rect 19165 18173 19199 18207
rect 20545 18173 20579 18207
rect 21005 18173 21039 18207
rect 21281 18173 21315 18207
rect 21649 18173 21683 18207
rect 21905 18173 21939 18207
rect 4629 18105 4663 18139
rect 11897 18105 11931 18139
rect 21557 18105 21591 18139
rect 5181 18037 5215 18071
rect 6561 18037 6595 18071
rect 7389 18037 7423 18071
rect 9781 18037 9815 18071
rect 15577 18037 15611 18071
rect 16681 18037 16715 18071
rect 16865 18037 16899 18071
rect 18705 18037 18739 18071
rect 21373 18037 21407 18071
rect 23029 18037 23063 18071
rect 5641 17833 5675 17867
rect 8677 17833 8711 17867
rect 10333 17833 10367 17867
rect 13093 17833 13127 17867
rect 16497 17833 16531 17867
rect 18153 17833 18187 17867
rect 21649 17833 21683 17867
rect 4629 17765 4663 17799
rect 4813 17765 4847 17799
rect 4997 17765 5031 17799
rect 5273 17765 5307 17799
rect 5825 17765 5859 17799
rect 7665 17765 7699 17799
rect 14013 17765 14047 17799
rect 16129 17765 16163 17799
rect 16345 17765 16379 17799
rect 18521 17765 18555 17799
rect 19042 17765 19076 17799
rect 23029 17765 23063 17799
rect 5089 17697 5123 17731
rect 5365 17697 5399 17731
rect 5457 17697 5491 17731
rect 6193 17697 6227 17731
rect 6837 17697 6871 17731
rect 8309 17697 8343 17731
rect 9965 17697 9999 17731
rect 10977 17697 11011 17731
rect 11161 17697 11195 17731
rect 12265 17697 12299 17731
rect 12725 17697 12759 17731
rect 13369 17697 13403 17731
rect 13829 17697 13863 17731
rect 15669 17697 15703 17731
rect 15761 17697 15795 17731
rect 15945 17697 15979 17731
rect 16773 17697 16807 17731
rect 17049 17697 17083 17731
rect 17233 17697 17267 17731
rect 17601 17697 17635 17731
rect 18061 17697 18095 17731
rect 18337 17697 18371 17731
rect 18429 17697 18463 17731
rect 18705 17697 18739 17731
rect 21833 17697 21867 17731
rect 21925 17697 21959 17731
rect 22385 17697 22419 17731
rect 22569 17697 22603 17731
rect 6009 17629 6043 17663
rect 6745 17629 6779 17663
rect 8217 17629 8251 17663
rect 10057 17629 10091 17663
rect 11069 17629 11103 17663
rect 11713 17629 11747 17663
rect 12357 17629 12391 17663
rect 12633 17629 12667 17663
rect 13277 17629 13311 17663
rect 17739 17629 17773 17663
rect 18797 17629 18831 17663
rect 21649 17629 21683 17663
rect 22293 17629 22327 17663
rect 6193 17561 6227 17595
rect 11989 17561 12023 17595
rect 16589 17561 16623 17595
rect 17877 17561 17911 17595
rect 13737 17493 13771 17527
rect 14197 17493 14231 17527
rect 16313 17493 16347 17527
rect 17969 17493 18003 17527
rect 20177 17493 20211 17527
rect 6285 17289 6319 17323
rect 11161 17289 11195 17323
rect 15025 17289 15059 17323
rect 16405 17289 16439 17323
rect 17141 17289 17175 17323
rect 17417 17289 17451 17323
rect 17693 17289 17727 17323
rect 18153 17289 18187 17323
rect 22385 17289 22419 17323
rect 6561 17221 6595 17255
rect 9229 17221 9263 17255
rect 14565 17221 14599 17255
rect 15485 17221 15519 17255
rect 16037 17221 16071 17255
rect 16957 17221 16991 17255
rect 17969 17221 18003 17255
rect 5089 17153 5123 17187
rect 10241 17153 10275 17187
rect 10701 17153 10735 17187
rect 15577 17153 15611 17187
rect 16313 17153 16347 17187
rect 17693 17153 17727 17187
rect 4905 17085 4939 17119
rect 5273 17085 5307 17119
rect 5365 17085 5399 17119
rect 5457 17085 5491 17119
rect 5615 17085 5649 17119
rect 5733 17085 5767 17119
rect 5917 17085 5951 17119
rect 6193 17085 6227 17119
rect 6377 17085 6411 17119
rect 6469 17085 6503 17119
rect 6837 17085 6871 17119
rect 7021 17085 7055 17119
rect 8861 17085 8895 17119
rect 8953 17085 8987 17119
rect 9413 17085 9447 17119
rect 9689 17085 9723 17119
rect 9873 17085 9907 17119
rect 10333 17085 10367 17119
rect 10793 17085 10827 17119
rect 14289 17085 14323 17119
rect 14565 17085 14599 17119
rect 14657 17085 14691 17119
rect 14841 17085 14875 17119
rect 15301 17085 15335 17119
rect 16589 17085 16623 17119
rect 16681 17085 16715 17119
rect 17049 17085 17083 17119
rect 17325 17085 17359 17119
rect 17601 17085 17635 17119
rect 18337 17085 18371 17119
rect 18521 17085 18555 17119
rect 18705 17085 18739 17119
rect 18961 17085 18995 17119
rect 20729 17085 20763 17119
rect 20821 17085 20855 17119
rect 22661 17085 22695 17119
rect 5825 17017 5859 17051
rect 6929 17017 6963 17051
rect 9137 17017 9171 17051
rect 15209 17017 15243 17051
rect 15669 17017 15703 17051
rect 16957 17017 16991 17051
rect 20545 17017 20579 17051
rect 21088 17017 21122 17051
rect 6101 16949 6135 16983
rect 9038 16949 9072 16983
rect 9965 16949 9999 16983
rect 14381 16949 14415 16983
rect 16773 16949 16807 16983
rect 20085 16949 20119 16983
rect 22201 16949 22235 16983
rect 5089 16745 5123 16779
rect 9505 16745 9539 16779
rect 10073 16745 10107 16779
rect 14473 16745 14507 16779
rect 19073 16745 19107 16779
rect 21281 16745 21315 16779
rect 9873 16677 9907 16711
rect 15945 16677 15979 16711
rect 4721 16609 4755 16643
rect 4905 16609 4939 16643
rect 6009 16609 6043 16643
rect 6837 16609 6871 16643
rect 7113 16609 7147 16643
rect 9321 16609 9355 16643
rect 9597 16609 9631 16643
rect 9781 16609 9815 16643
rect 14657 16609 14691 16643
rect 14841 16609 14875 16643
rect 14933 16609 14967 16643
rect 15025 16609 15059 16643
rect 15209 16609 15243 16643
rect 15669 16609 15703 16643
rect 16313 16609 16347 16643
rect 16589 16609 16623 16643
rect 16957 16609 16991 16643
rect 17049 16609 17083 16643
rect 17141 16609 17175 16643
rect 18429 16609 18463 16643
rect 18613 16609 18647 16643
rect 19073 16609 19107 16643
rect 19257 16609 19291 16643
rect 21465 16609 21499 16643
rect 21649 16609 21683 16643
rect 21741 16609 21775 16643
rect 6101 16541 6135 16575
rect 6745 16541 6779 16575
rect 15117 16541 15151 16575
rect 15761 16541 15795 16575
rect 15945 16541 15979 16575
rect 16405 16541 16439 16575
rect 16865 16541 16899 16575
rect 6469 16473 6503 16507
rect 7389 16473 7423 16507
rect 16497 16473 16531 16507
rect 18429 16473 18463 16507
rect 6377 16405 6411 16439
rect 7573 16405 7607 16439
rect 10057 16405 10091 16439
rect 10241 16405 10275 16439
rect 16129 16405 16163 16439
rect 17325 16405 17359 16439
rect 7573 16201 7607 16235
rect 15301 16201 15335 16235
rect 15485 16201 15519 16235
rect 17233 16201 17267 16235
rect 19441 16201 19475 16235
rect 21373 16201 21407 16235
rect 21833 16201 21867 16235
rect 5181 16133 5215 16167
rect 6837 16133 6871 16167
rect 8953 16133 8987 16167
rect 13829 16133 13863 16167
rect 19993 16133 20027 16167
rect 6561 16065 6595 16099
rect 6929 16065 6963 16099
rect 7389 16065 7423 16099
rect 7757 16065 7791 16099
rect 8493 16065 8527 16099
rect 9413 16065 9447 16099
rect 11805 16065 11839 16099
rect 12265 16065 12299 16099
rect 12633 16065 12667 16099
rect 14565 16065 14599 16099
rect 19809 16065 19843 16099
rect 21557 16065 21591 16099
rect 4905 15997 4939 16031
rect 6469 15997 6503 16031
rect 7297 15997 7331 16031
rect 7849 15997 7883 16031
rect 8585 15997 8619 16031
rect 9505 15997 9539 16031
rect 10793 15997 10827 16031
rect 10886 15997 10920 16031
rect 11897 15997 11931 16031
rect 12541 15997 12575 16031
rect 13001 15997 13035 16031
rect 13185 15997 13219 16031
rect 13553 15997 13587 16031
rect 14657 15997 14691 16031
rect 14933 15997 14967 16031
rect 15393 15997 15427 16031
rect 15577 15997 15611 16031
rect 16129 15997 16163 16031
rect 16313 15997 16347 16031
rect 16497 15997 16531 16031
rect 16957 15997 16991 16031
rect 17049 15997 17083 16031
rect 17325 15997 17359 16031
rect 19349 15997 19383 16031
rect 19533 15997 19567 16031
rect 20085 15997 20119 16031
rect 20545 15997 20579 16031
rect 20821 15997 20855 16031
rect 21005 15997 21039 16031
rect 21281 15997 21315 16031
rect 21649 15997 21683 16031
rect 21741 15997 21775 16031
rect 22385 15997 22419 16031
rect 4997 15929 5031 15963
rect 5181 15929 5215 15963
rect 13369 15929 13403 15963
rect 13829 15929 13863 15963
rect 15117 15929 15151 15963
rect 16405 15929 16439 15963
rect 20729 15929 20763 15963
rect 21557 15929 21591 15963
rect 22201 15929 22235 15963
rect 8217 15861 8251 15895
rect 9873 15861 9907 15895
rect 11161 15861 11195 15895
rect 12909 15861 12943 15895
rect 13645 15861 13679 15895
rect 14289 15861 14323 15895
rect 16681 15861 16715 15895
rect 16773 15861 16807 15895
rect 19717 15861 19751 15895
rect 19809 15861 19843 15895
rect 20361 15861 20395 15895
rect 20913 15861 20947 15895
rect 22017 15861 22051 15895
rect 22569 15861 22603 15895
rect 5641 15657 5675 15691
rect 7573 15657 7607 15691
rect 8493 15657 8527 15691
rect 17509 15657 17543 15691
rect 20295 15657 20329 15691
rect 5273 15589 5307 15623
rect 6070 15589 6104 15623
rect 7757 15589 7791 15623
rect 16396 15589 16430 15623
rect 20085 15589 20119 15623
rect 5089 15521 5123 15555
rect 5365 15521 5399 15555
rect 5457 15521 5491 15555
rect 7481 15521 7515 15555
rect 8125 15521 8159 15555
rect 8585 15521 8619 15555
rect 8678 15521 8712 15555
rect 9597 15521 9631 15555
rect 9690 15521 9724 15555
rect 10517 15521 10551 15555
rect 11253 15521 11287 15555
rect 11713 15521 11747 15555
rect 11897 15521 11931 15555
rect 11989 15521 12023 15555
rect 12081 15521 12115 15555
rect 12265 15521 12299 15555
rect 12541 15521 12575 15555
rect 12633 15521 12667 15555
rect 12817 15521 12851 15555
rect 14565 15521 14599 15555
rect 14749 15521 14783 15555
rect 17693 15521 17727 15555
rect 17877 15521 17911 15555
rect 18797 15521 18831 15555
rect 19717 15521 19751 15555
rect 19901 15521 19935 15555
rect 20545 15521 20579 15555
rect 20821 15521 20855 15555
rect 21649 15521 21683 15555
rect 22293 15521 22327 15555
rect 5825 15453 5859 15487
rect 8033 15453 8067 15487
rect 9965 15453 9999 15487
rect 10425 15453 10459 15487
rect 11161 15453 11195 15487
rect 12173 15453 12207 15487
rect 13829 15453 13863 15487
rect 16129 15453 16163 15487
rect 18889 15453 18923 15487
rect 20637 15453 20671 15487
rect 21557 15453 21591 15487
rect 22201 15453 22235 15487
rect 7757 15385 7791 15419
rect 10149 15385 10183 15419
rect 20453 15385 20487 15419
rect 21005 15385 21039 15419
rect 7205 15317 7239 15351
rect 8769 15317 8803 15351
rect 11529 15317 11563 15351
rect 11713 15317 11747 15351
rect 13001 15317 13035 15351
rect 17785 15317 17819 15351
rect 18429 15317 18463 15351
rect 19809 15317 19843 15351
rect 20269 15317 20303 15351
rect 20637 15317 20671 15351
rect 21281 15317 21315 15351
rect 21925 15317 21959 15351
rect 10977 15113 11011 15147
rect 12173 15113 12207 15147
rect 12909 15113 12943 15147
rect 13921 15113 13955 15147
rect 14933 15113 14967 15147
rect 17877 15113 17911 15147
rect 18337 15113 18371 15147
rect 20729 15113 20763 15147
rect 13093 15045 13127 15079
rect 14289 15045 14323 15079
rect 21833 15045 21867 15079
rect 22109 15045 22143 15079
rect 8953 14977 8987 15011
rect 9229 14977 9263 15011
rect 13829 14977 13863 15011
rect 19809 14977 19843 15011
rect 20269 14977 20303 15011
rect 21373 14977 21407 15011
rect 21925 14977 21959 15011
rect 22477 14977 22511 15011
rect 8861 14909 8895 14943
rect 9321 14909 9355 14943
rect 9414 14909 9448 14943
rect 9873 14909 9907 14943
rect 10057 14909 10091 14943
rect 10425 14909 10459 14943
rect 11437 14909 11471 14943
rect 11713 14909 11747 14943
rect 13553 14909 13587 14943
rect 14013 14909 14047 14943
rect 14381 14909 14415 14943
rect 14473 14909 14507 14943
rect 14657 14909 14691 14943
rect 14749 14909 14783 14943
rect 16497 14909 16531 14943
rect 16764 14909 16798 14943
rect 18153 14909 18187 14943
rect 19901 14909 19935 14943
rect 20453 14909 20487 14943
rect 21465 14909 21499 14943
rect 22017 14909 22051 14943
rect 22385 14909 22419 14943
rect 22661 14909 22695 14943
rect 22753 14909 22787 14943
rect 10241 14841 10275 14875
rect 10793 14841 10827 14875
rect 11989 14841 12023 14875
rect 12189 14841 12223 14875
rect 12725 14841 12759 14875
rect 12925 14841 12959 14875
rect 17969 14841 18003 14875
rect 18705 14841 18739 14875
rect 18889 14841 18923 14875
rect 20545 14841 20579 14875
rect 20729 14841 20763 14875
rect 22293 14841 22327 14875
rect 9689 14773 9723 14807
rect 10057 14773 10091 14807
rect 10609 14773 10643 14807
rect 10993 14773 11027 14807
rect 11161 14773 11195 14807
rect 11529 14773 11563 14807
rect 11897 14773 11931 14807
rect 12357 14773 12391 14807
rect 13645 14773 13679 14807
rect 19073 14773 19107 14807
rect 22477 14773 22511 14807
rect 6193 14569 6227 14603
rect 10609 14569 10643 14603
rect 12909 14569 12943 14603
rect 14539 14569 14573 14603
rect 15025 14569 15059 14603
rect 17515 14569 17549 14603
rect 19073 14569 19107 14603
rect 22201 14569 22235 14603
rect 9689 14501 9723 14535
rect 9873 14501 9907 14535
rect 11253 14501 11287 14535
rect 11345 14501 11379 14535
rect 13921 14501 13955 14535
rect 14749 14501 14783 14535
rect 14841 14501 14875 14535
rect 17601 14501 17635 14535
rect 19225 14501 19259 14535
rect 19441 14501 19475 14535
rect 22569 14501 22603 14535
rect 22661 14501 22695 14535
rect 6285 14433 6319 14467
rect 9229 14433 9263 14467
rect 9413 14433 9447 14467
rect 9965 14433 9999 14467
rect 10241 14433 10275 14467
rect 10425 14433 10459 14467
rect 11161 14433 11195 14467
rect 11529 14433 11563 14467
rect 11621 14433 11655 14467
rect 11897 14433 11931 14467
rect 11989 14433 12023 14467
rect 12817 14433 12851 14467
rect 13093 14433 13127 14467
rect 13369 14433 13403 14467
rect 13553 14433 13587 14467
rect 13829 14433 13863 14467
rect 14105 14433 14139 14467
rect 15117 14433 15151 14467
rect 16681 14433 16715 14467
rect 17417 14433 17451 14467
rect 17693 14433 17727 14467
rect 17785 14433 17819 14467
rect 17969 14433 18003 14467
rect 18613 14433 18647 14467
rect 21557 14433 21591 14467
rect 22017 14433 22051 14467
rect 22293 14433 22327 14467
rect 22477 14433 22511 14467
rect 22779 14433 22813 14467
rect 6377 14365 6411 14399
rect 11713 14365 11747 14399
rect 13277 14365 13311 14399
rect 16957 14365 16991 14399
rect 18153 14365 18187 14399
rect 18521 14365 18555 14399
rect 21925 14365 21959 14399
rect 22937 14365 22971 14399
rect 9413 14297 9447 14331
rect 10977 14297 11011 14331
rect 16865 14297 16899 14331
rect 5825 14229 5859 14263
rect 9505 14229 9539 14263
rect 10149 14229 10183 14263
rect 11805 14229 11839 14263
rect 13461 14229 13495 14263
rect 14289 14229 14323 14263
rect 14381 14229 14415 14263
rect 14565 14229 14599 14263
rect 14841 14229 14875 14263
rect 16773 14229 16807 14263
rect 18889 14229 18923 14263
rect 19257 14229 19291 14263
rect 22017 14229 22051 14263
rect 4261 14025 4295 14059
rect 8953 14025 8987 14059
rect 10977 14025 11011 14059
rect 14657 14025 14691 14059
rect 16957 14025 16991 14059
rect 17325 14025 17359 14059
rect 17785 14025 17819 14059
rect 17969 14025 18003 14059
rect 18061 14025 18095 14059
rect 19073 14025 19107 14059
rect 19257 14025 19291 14059
rect 21741 14025 21775 14059
rect 21925 14025 21959 14059
rect 5733 13957 5767 13991
rect 7205 13957 7239 13991
rect 14749 13957 14783 13991
rect 7665 13889 7699 13923
rect 7849 13889 7883 13923
rect 10793 13889 10827 13923
rect 13093 13889 13127 13923
rect 13185 13889 13219 13923
rect 13277 13889 13311 13923
rect 14841 13889 14875 13923
rect 18889 13889 18923 13923
rect 20361 13889 20395 13923
rect 5385 13821 5419 13855
rect 5641 13821 5675 13855
rect 6857 13821 6891 13855
rect 7113 13821 7147 13855
rect 8953 13821 8987 13855
rect 9137 13821 9171 13855
rect 9229 13821 9263 13855
rect 9781 13821 9815 13855
rect 9965 13821 9999 13855
rect 10057 13821 10091 13855
rect 10241 13821 10275 13855
rect 10609 13821 10643 13855
rect 10885 13821 10919 13855
rect 11069 13821 11103 13855
rect 13001 13821 13035 13855
rect 13737 13821 13771 13855
rect 13891 13821 13925 13855
rect 14565 13821 14599 13855
rect 15485 13821 15519 13855
rect 16957 13821 16991 13855
rect 17049 13821 17083 13855
rect 18061 13821 18095 13855
rect 18337 13821 18371 13855
rect 18797 13821 18831 13855
rect 19073 13821 19107 13855
rect 20085 13821 20119 13855
rect 20269 13821 20303 13855
rect 20628 13821 20662 13855
rect 22109 13821 22143 13855
rect 22201 13821 22235 13855
rect 7573 13753 7607 13787
rect 15752 13753 15786 13787
rect 17601 13753 17635 13787
rect 17817 13753 17851 13787
rect 21925 13753 21959 13787
rect 9597 13685 9631 13719
rect 10149 13685 10183 13719
rect 10425 13685 10459 13719
rect 12817 13685 12851 13719
rect 14105 13685 14139 13719
rect 16865 13685 16899 13719
rect 18245 13685 18279 13719
rect 19901 13685 19935 13719
rect 5825 13481 5859 13515
rect 6193 13481 6227 13515
rect 12449 13481 12483 13515
rect 16129 13481 16163 13515
rect 18537 13481 18571 13515
rect 6285 13413 6319 13447
rect 16497 13413 16531 13447
rect 18337 13413 18371 13447
rect 19901 13413 19935 13447
rect 21281 13413 21315 13447
rect 21481 13413 21515 13447
rect 21741 13413 21775 13447
rect 21941 13413 21975 13447
rect 7021 13345 7055 13379
rect 7288 13345 7322 13379
rect 8769 13345 8803 13379
rect 8953 13345 8987 13379
rect 9229 13345 9263 13379
rect 9321 13345 9355 13379
rect 9413 13345 9447 13379
rect 9597 13345 9631 13379
rect 9965 13345 9999 13379
rect 10241 13345 10275 13379
rect 11805 13345 11839 13379
rect 11897 13345 11931 13379
rect 12357 13345 12391 13379
rect 12817 13345 12851 13379
rect 12909 13345 12943 13379
rect 14289 13345 14323 13379
rect 14381 13345 14415 13379
rect 14473 13345 14507 13379
rect 14933 13345 14967 13379
rect 20269 13345 20303 13379
rect 22385 13345 22419 13379
rect 22569 13345 22603 13379
rect 22845 13345 22879 13379
rect 6469 13277 6503 13311
rect 9689 13277 9723 13311
rect 10333 13277 10367 13311
rect 11989 13277 12023 13311
rect 12081 13277 12115 13311
rect 14565 13277 14599 13311
rect 14749 13277 14783 13311
rect 15117 13277 15151 13311
rect 16589 13277 16623 13311
rect 16773 13277 16807 13311
rect 20453 13277 20487 13311
rect 20545 13277 20579 13311
rect 20637 13277 20671 13311
rect 20729 13277 20763 13311
rect 22201 13277 22235 13311
rect 8861 13209 8895 13243
rect 9781 13209 9815 13243
rect 18705 13209 18739 13243
rect 22661 13209 22695 13243
rect 8401 13141 8435 13175
rect 9045 13141 9079 13175
rect 10149 13141 10183 13175
rect 11621 13141 11655 13175
rect 12725 13141 12759 13175
rect 14105 13141 14139 13175
rect 18521 13141 18555 13175
rect 19717 13141 19751 13175
rect 19901 13141 19935 13175
rect 20913 13141 20947 13175
rect 21465 13141 21499 13175
rect 21649 13141 21683 13175
rect 21925 13141 21959 13175
rect 22109 13141 22143 13175
rect 6561 12937 6595 12971
rect 7481 12937 7515 12971
rect 11897 12937 11931 12971
rect 15301 12937 15335 12971
rect 18153 12937 18187 12971
rect 18705 12937 18739 12971
rect 21005 12937 21039 12971
rect 21097 12937 21131 12971
rect 21281 12937 21315 12971
rect 21925 12937 21959 12971
rect 22753 12937 22787 12971
rect 18521 12869 18555 12903
rect 22845 12869 22879 12903
rect 6285 12801 6319 12835
rect 8125 12801 8159 12835
rect 10333 12801 10367 12835
rect 15853 12801 15887 12835
rect 16037 12801 16071 12835
rect 6018 12733 6052 12767
rect 6377 12733 6411 12767
rect 6561 12733 6595 12767
rect 7849 12733 7883 12767
rect 8585 12733 8619 12767
rect 10425 12733 10459 12767
rect 11621 12733 11655 12767
rect 11713 12733 11747 12767
rect 13102 12733 13136 12767
rect 13369 12733 13403 12767
rect 13921 12733 13955 12767
rect 14188 12733 14222 12767
rect 17693 12733 17727 12767
rect 17877 12733 17911 12767
rect 18889 12733 18923 12767
rect 19165 12733 19199 12767
rect 19625 12733 19659 12767
rect 19881 12733 19915 12767
rect 21649 12733 21683 12767
rect 22293 12733 22327 12767
rect 23029 12733 23063 12767
rect 7941 12665 7975 12699
rect 8852 12665 8886 12699
rect 17785 12665 17819 12699
rect 19073 12665 19107 12699
rect 19257 12665 19291 12699
rect 19441 12665 19475 12699
rect 21281 12665 21315 12699
rect 22385 12665 22419 12699
rect 22569 12665 22603 12699
rect 4905 12597 4939 12631
rect 6745 12597 6779 12631
rect 9965 12597 9999 12631
rect 10793 12597 10827 12631
rect 11989 12597 12023 12631
rect 15393 12597 15427 12631
rect 15761 12597 15795 12631
rect 17969 12597 18003 12631
rect 18153 12597 18187 12631
rect 21741 12597 21775 12631
rect 21925 12597 21959 12631
rect 5641 12393 5675 12427
rect 12725 12393 12759 12427
rect 13553 12393 13587 12427
rect 19073 12393 19107 12427
rect 20637 12393 20671 12427
rect 6469 12325 6503 12359
rect 11612 12325 11646 12359
rect 17417 12325 17451 12359
rect 17960 12325 17994 12359
rect 21894 12325 21928 12359
rect 5365 12257 5399 12291
rect 5457 12257 5491 12291
rect 6193 12257 6227 12291
rect 6745 12257 6779 12291
rect 7113 12257 7147 12291
rect 7297 12257 7331 12291
rect 9229 12257 9263 12291
rect 13737 12257 13771 12291
rect 13921 12257 13955 12291
rect 14361 12257 14395 12291
rect 16497 12257 16531 12291
rect 17601 12257 17635 12291
rect 19421 12257 19455 12291
rect 20821 12257 20855 12291
rect 21005 12257 21039 12291
rect 21373 12257 21407 12291
rect 5641 12189 5675 12223
rect 6285 12189 6319 12223
rect 6561 12189 6595 12223
rect 9321 12189 9355 12223
rect 11345 12189 11379 12223
rect 14013 12189 14047 12223
rect 14105 12189 14139 12223
rect 16589 12189 16623 12223
rect 17693 12189 17727 12223
rect 19165 12189 19199 12223
rect 21649 12189 21683 12223
rect 6929 12121 6963 12155
rect 5825 12053 5859 12087
rect 6469 12053 6503 12087
rect 7205 12053 7239 12087
rect 9505 12053 9539 12087
rect 15485 12053 15519 12087
rect 16865 12053 16899 12087
rect 17233 12053 17267 12087
rect 20545 12053 20579 12087
rect 21465 12053 21499 12087
rect 23029 12053 23063 12087
rect 6653 11849 6687 11883
rect 16037 11849 16071 11883
rect 16129 11849 16163 11883
rect 16589 11849 16623 11883
rect 17049 11849 17083 11883
rect 18061 11849 18095 11883
rect 18245 11849 18279 11883
rect 19441 11849 19475 11883
rect 21097 11849 21131 11883
rect 21557 11849 21591 11883
rect 6929 11781 6963 11815
rect 17509 11781 17543 11815
rect 5917 11713 5951 11747
rect 8585 11713 8619 11747
rect 8769 11713 8803 11747
rect 16221 11713 16255 11747
rect 21189 11713 21223 11747
rect 6009 11645 6043 11679
rect 7113 11645 7147 11679
rect 7205 11645 7239 11679
rect 8493 11645 8527 11679
rect 8861 11645 8895 11679
rect 10977 11645 11011 11679
rect 14657 11645 14691 11679
rect 14924 11645 14958 11679
rect 16405 11645 16439 11679
rect 17233 11645 17267 11679
rect 17325 11645 17359 11679
rect 19717 11645 19751 11679
rect 21373 11645 21407 11679
rect 21649 11645 21683 11679
rect 6469 11577 6503 11611
rect 6929 11577 6963 11611
rect 9128 11577 9162 11611
rect 11244 11577 11278 11611
rect 16129 11577 16163 11611
rect 17049 11577 17083 11611
rect 17877 11577 17911 11611
rect 18077 11577 18111 11611
rect 19257 11577 19291 11611
rect 19962 11577 19996 11611
rect 21894 11577 21928 11611
rect 6377 11509 6411 11543
rect 6669 11509 6703 11543
rect 6837 11509 6871 11543
rect 8769 11509 8803 11543
rect 10241 11509 10275 11543
rect 12357 11509 12391 11543
rect 19457 11509 19491 11543
rect 19625 11509 19659 11543
rect 23029 11509 23063 11543
rect 5483 11305 5517 11339
rect 7113 11305 7147 11339
rect 7481 11305 7515 11339
rect 8125 11305 8159 11339
rect 9413 11305 9447 11339
rect 9873 11305 9907 11339
rect 10701 11305 10735 11339
rect 11253 11305 11287 11339
rect 11713 11305 11747 11339
rect 15485 11305 15519 11339
rect 16605 11305 16639 11339
rect 16773 11305 16807 11339
rect 17417 11305 17451 11339
rect 17785 11305 17819 11339
rect 18061 11305 18095 11339
rect 20085 11305 20119 11339
rect 20545 11305 20579 11339
rect 21557 11305 21591 11339
rect 21741 11305 21775 11339
rect 5273 11237 5307 11271
rect 6193 11237 6227 11271
rect 6377 11237 6411 11271
rect 8369 11237 8403 11271
rect 8585 11237 8619 11271
rect 15945 11237 15979 11271
rect 16405 11237 16439 11271
rect 17509 11237 17543 11271
rect 18337 11237 18371 11271
rect 20453 11237 20487 11271
rect 22569 11237 22603 11271
rect 4997 11169 5031 11203
rect 5181 11169 5215 11203
rect 5825 11169 5859 11203
rect 6009 11169 6043 11203
rect 6285 11169 6319 11203
rect 6653 11169 6687 11203
rect 6837 11169 6871 11203
rect 7113 11169 7147 11203
rect 7297 11169 7331 11203
rect 7389 11169 7423 11203
rect 7665 11169 7699 11203
rect 7757 11169 7791 11203
rect 8953 11169 8987 11203
rect 9781 11169 9815 11203
rect 10241 11169 10275 11203
rect 10517 11169 10551 11203
rect 10977 11169 11011 11203
rect 11161 11169 11195 11203
rect 11621 11169 11655 11203
rect 12265 11169 12299 11203
rect 12541 11169 12575 11203
rect 12725 11169 12759 11203
rect 12817 11169 12851 11203
rect 14289 11169 14323 11203
rect 14473 11169 14507 11203
rect 14749 11169 14783 11203
rect 15025 11169 15059 11203
rect 15301 11169 15335 11203
rect 15485 11169 15519 11203
rect 15669 11169 15703 11203
rect 15761 11169 15795 11203
rect 17049 11169 17083 11203
rect 17693 11169 17727 11203
rect 17877 11169 17911 11203
rect 18705 11169 18739 11203
rect 20269 11169 20303 11203
rect 20545 11169 20579 11203
rect 20729 11169 20763 11203
rect 22109 11169 22143 11203
rect 22385 11169 22419 11203
rect 7849 11101 7883 11135
rect 9045 11101 9079 11135
rect 9965 11101 9999 11135
rect 10333 11101 10367 11135
rect 11069 11101 11103 11135
rect 11805 11101 11839 11135
rect 12449 11101 12483 11135
rect 14565 11101 14599 11135
rect 16957 11101 16991 11135
rect 7021 11033 7055 11067
rect 8217 11033 8251 11067
rect 13001 11033 13035 11067
rect 15163 11033 15197 11067
rect 15945 11033 15979 11067
rect 4813 10965 4847 10999
rect 5457 10965 5491 10999
rect 5641 10965 5675 10999
rect 6837 10965 6871 10999
rect 7665 10965 7699 10999
rect 7757 10965 7791 10999
rect 8401 10965 8435 10999
rect 9137 10965 9171 10999
rect 9321 10965 9355 10999
rect 10241 10965 10275 10999
rect 12081 10965 12115 10999
rect 12633 10965 12667 10999
rect 14289 10965 14323 10999
rect 14933 10965 14967 10999
rect 16589 10965 16623 10999
rect 18153 10965 18187 10999
rect 18337 10965 18371 10999
rect 21741 10965 21775 10999
rect 22201 10965 22235 10999
rect 6285 10761 6319 10795
rect 9505 10761 9539 10795
rect 12541 10761 12575 10795
rect 17049 10761 17083 10795
rect 21465 10761 21499 10795
rect 22385 10761 22419 10795
rect 22753 10761 22787 10795
rect 10425 10693 10459 10727
rect 12403 10693 12437 10727
rect 17141 10693 17175 10727
rect 8493 10625 8527 10659
rect 8953 10625 8987 10659
rect 9873 10625 9907 10659
rect 11713 10625 11747 10659
rect 14565 10625 14599 10659
rect 22293 10625 22327 10659
rect 4629 10557 4663 10591
rect 4813 10557 4847 10591
rect 4905 10557 4939 10591
rect 6561 10557 6595 10591
rect 8585 10557 8619 10591
rect 9965 10557 9999 10591
rect 10425 10557 10459 10591
rect 10609 10557 10643 10591
rect 10701 10557 10735 10591
rect 11345 10557 11379 10591
rect 11529 10557 11563 10591
rect 11805 10557 11839 10591
rect 12265 10557 12299 10591
rect 12725 10557 12759 10591
rect 13553 10557 13587 10591
rect 13737 10557 13771 10591
rect 14657 10557 14691 10591
rect 15117 10557 15151 10591
rect 15301 10557 15335 10591
rect 16865 10557 16899 10591
rect 18254 10557 18288 10591
rect 18521 10557 18555 10591
rect 20821 10557 20855 10591
rect 21833 10557 21867 10591
rect 22109 10557 22143 10591
rect 22385 10557 22419 10591
rect 22569 10557 22603 10591
rect 5172 10489 5206 10523
rect 6377 10489 6411 10523
rect 9321 10489 9355 10523
rect 12633 10489 12667 10523
rect 15209 10489 15243 10523
rect 16681 10489 16715 10523
rect 21005 10489 21039 10523
rect 21189 10489 21223 10523
rect 21465 10489 21499 10523
rect 4721 10421 4755 10455
rect 6745 10421 6779 10455
rect 9521 10421 9555 10455
rect 9689 10421 9723 10455
rect 10333 10421 10367 10455
rect 11437 10421 11471 10455
rect 12173 10421 12207 10455
rect 13737 10421 13771 10455
rect 15025 10421 15059 10455
rect 21281 10421 21315 10455
rect 21925 10421 21959 10455
rect 4353 10217 4387 10251
rect 9873 10217 9907 10251
rect 16405 10217 16439 10251
rect 16865 10217 16899 10251
rect 21281 10217 21315 10251
rect 22109 10217 22143 10251
rect 3985 10149 4019 10183
rect 4813 10149 4847 10183
rect 5089 10149 5123 10183
rect 5365 10149 5399 10183
rect 9413 10149 9447 10183
rect 12173 10149 12207 10183
rect 21097 10149 21131 10183
rect 22569 10149 22603 10183
rect 4215 10115 4249 10149
rect 4445 10081 4479 10115
rect 5273 10081 5307 10115
rect 5457 10081 5491 10115
rect 6938 10081 6972 10115
rect 7205 10081 7239 10115
rect 8769 10081 8803 10115
rect 9689 10081 9723 10115
rect 11713 10081 11747 10115
rect 12449 10081 12483 10115
rect 13829 10081 13863 10115
rect 14565 10081 14599 10115
rect 15209 10081 15243 10115
rect 16313 10081 16347 10115
rect 16589 10081 16623 10115
rect 17978 10081 18012 10115
rect 18245 10081 18279 10115
rect 19717 10081 19751 10115
rect 20729 10081 20763 10115
rect 20821 10081 20855 10115
rect 20913 10081 20947 10115
rect 21649 10081 21683 10115
rect 22477 10081 22511 10115
rect 22753 10081 22787 10115
rect 8861 10013 8895 10047
rect 9505 10013 9539 10047
rect 11621 10013 11655 10047
rect 12265 10013 12299 10047
rect 13737 10013 13771 10047
rect 14657 10013 14691 10047
rect 15117 10013 15151 10047
rect 19901 10013 19935 10047
rect 20545 10013 20579 10047
rect 21465 10013 21499 10047
rect 21557 10013 21591 10047
rect 21741 10013 21775 10047
rect 9137 9945 9171 9979
rect 14197 9945 14231 9979
rect 4169 9877 4203 9911
rect 4813 9877 4847 9911
rect 4997 9877 5031 9911
rect 5641 9877 5675 9911
rect 5825 9877 5859 9911
rect 9689 9877 9723 9911
rect 11989 9877 12023 9911
rect 12173 9877 12207 9911
rect 12633 9877 12667 9911
rect 14841 9877 14875 9911
rect 15485 9877 15519 9911
rect 16773 9877 16807 9911
rect 19533 9877 19567 9911
rect 21925 9877 21959 9911
rect 22109 9877 22143 9911
rect 22937 9877 22971 9911
rect 4629 9673 4663 9707
rect 4813 9673 4847 9707
rect 6745 9673 6779 9707
rect 6929 9673 6963 9707
rect 8769 9673 8803 9707
rect 11345 9673 11379 9707
rect 14381 9673 14415 9707
rect 15025 9673 15059 9707
rect 17325 9673 17359 9707
rect 17601 9673 17635 9707
rect 17785 9673 17819 9707
rect 19257 9673 19291 9707
rect 21189 9673 21223 9707
rect 6285 9605 6319 9639
rect 12449 9605 12483 9639
rect 14565 9605 14599 9639
rect 15485 9605 15519 9639
rect 16957 9605 16991 9639
rect 17509 9605 17543 9639
rect 4905 9537 4939 9571
rect 10885 9537 10919 9571
rect 12173 9537 12207 9571
rect 15209 9537 15243 9571
rect 5161 9469 5195 9503
rect 6377 9469 6411 9503
rect 7941 9469 7975 9503
rect 8401 9469 8435 9503
rect 9045 9469 9079 9503
rect 9229 9469 9263 9503
rect 10977 9469 11011 9503
rect 12081 9469 12115 9503
rect 15025 9469 15059 9503
rect 15301 9469 15335 9503
rect 16681 9469 16715 9503
rect 16865 9469 16899 9503
rect 18797 9469 18831 9503
rect 18981 9469 19015 9503
rect 19625 9469 19659 9503
rect 19809 9469 19843 9503
rect 21557 9469 21591 9503
rect 21824 9469 21858 9503
rect 4445 9401 4479 9435
rect 4661 9401 4695 9435
rect 6745 9401 6779 9435
rect 7757 9401 7791 9435
rect 14197 9401 14231 9435
rect 14413 9401 14447 9435
rect 17769 9401 17803 9435
rect 17969 9401 18003 9435
rect 20076 9401 20110 9435
rect 7573 9333 7607 9367
rect 8769 9333 8803 9367
rect 8953 9333 8987 9367
rect 9413 9333 9447 9367
rect 16865 9333 16899 9367
rect 17325 9333 17359 9367
rect 18797 9333 18831 9367
rect 19073 9333 19107 9367
rect 19257 9333 19291 9367
rect 22937 9333 22971 9367
rect 5273 9129 5307 9163
rect 7139 9129 7173 9163
rect 9137 9129 9171 9163
rect 9965 9129 9999 9163
rect 11145 9129 11179 9163
rect 11805 9129 11839 9163
rect 18455 9129 18489 9163
rect 20177 9129 20211 9163
rect 22753 9129 22787 9163
rect 5457 9061 5491 9095
rect 6929 9061 6963 9095
rect 9045 9061 9079 9095
rect 10609 9061 10643 9095
rect 11345 9061 11379 9095
rect 11713 9061 11747 9095
rect 13093 9061 13127 9095
rect 13277 9061 13311 9095
rect 14105 9061 14139 9095
rect 15209 9061 15243 9095
rect 15393 9061 15427 9095
rect 18245 9061 18279 9095
rect 20361 9061 20395 9095
rect 20913 9061 20947 9095
rect 21618 9061 21652 9095
rect 5641 8993 5675 9027
rect 7645 8993 7679 9027
rect 9229 8993 9263 9027
rect 9505 8993 9539 9027
rect 9597 8993 9631 9027
rect 9781 8993 9815 9027
rect 10149 8993 10183 9027
rect 10333 8993 10367 9027
rect 10793 8993 10827 9027
rect 11437 8993 11471 9027
rect 11621 8993 11655 9027
rect 12081 8993 12115 9027
rect 12265 8993 12299 9027
rect 13645 8993 13679 9027
rect 13829 8993 13863 9027
rect 14473 8993 14507 9027
rect 14749 8993 14783 9027
rect 14841 8993 14875 9027
rect 14933 8993 14967 9027
rect 16129 8993 16163 9027
rect 16313 8993 16347 9027
rect 17610 8993 17644 9027
rect 17877 8993 17911 9027
rect 18961 8993 18995 9027
rect 20729 8993 20763 9027
rect 7389 8925 7423 8959
rect 9413 8925 9447 8959
rect 18705 8925 18739 8959
rect 21097 8925 21131 8959
rect 21373 8925 21407 8959
rect 7297 8857 7331 8891
rect 8769 8857 8803 8891
rect 8861 8857 8895 8891
rect 10977 8857 11011 8891
rect 14565 8857 14599 8891
rect 15117 8857 15151 8891
rect 16497 8857 16531 8891
rect 18613 8857 18647 8891
rect 20085 8857 20119 8891
rect 7113 8789 7147 8823
rect 10241 8789 10275 8823
rect 10425 8789 10459 8823
rect 11161 8789 11195 8823
rect 11989 8789 12023 8823
rect 12449 8789 12483 8823
rect 13461 8789 13495 8823
rect 13921 8789 13955 8823
rect 14105 8789 14139 8823
rect 15577 8789 15611 8823
rect 18429 8789 18463 8823
rect 20361 8789 20395 8823
rect 7665 8585 7699 8619
rect 8033 8585 8067 8619
rect 8217 8585 8251 8619
rect 9965 8585 9999 8619
rect 10333 8585 10367 8619
rect 11161 8585 11195 8619
rect 12817 8585 12851 8619
rect 13185 8585 13219 8619
rect 13645 8585 13679 8619
rect 15301 8585 15335 8619
rect 17417 8585 17451 8619
rect 17601 8585 17635 8619
rect 20453 8585 20487 8619
rect 21741 8585 21775 8619
rect 22201 8585 22235 8619
rect 22477 8585 22511 8619
rect 10149 8517 10183 8551
rect 11345 8517 11379 8551
rect 20269 8517 20303 8551
rect 22293 8517 22327 8551
rect 22753 8517 22787 8551
rect 10701 8449 10735 8483
rect 10793 8449 10827 8483
rect 18889 8449 18923 8483
rect 21649 8449 21683 8483
rect 21833 8449 21867 8483
rect 5917 8381 5951 8415
rect 7573 8381 7607 8415
rect 7757 8381 7791 8415
rect 8585 8381 8619 8415
rect 11437 8381 11471 8415
rect 11693 8381 11727 8415
rect 13553 8381 13587 8415
rect 13737 8381 13771 8415
rect 13829 8381 13863 8415
rect 14085 8381 14119 8415
rect 16681 8381 16715 8415
rect 16957 8381 16991 8415
rect 17141 8381 17175 8415
rect 19156 8381 19190 8415
rect 20637 8381 20671 8415
rect 20897 8381 20931 8415
rect 21005 8381 21039 8415
rect 21189 8381 21223 8415
rect 21281 8381 21315 8415
rect 21373 8381 21407 8415
rect 22017 8381 22051 8415
rect 22937 8381 22971 8415
rect 5733 8313 5767 8347
rect 6101 8313 6135 8347
rect 7849 8313 7883 8347
rect 8852 8313 8886 8347
rect 10333 8313 10367 8347
rect 11161 8313 11195 8347
rect 13001 8313 13035 8347
rect 13217 8313 13251 8347
rect 16414 8313 16448 8347
rect 16773 8313 16807 8347
rect 17233 8313 17267 8347
rect 17433 8313 17467 8347
rect 21741 8313 21775 8347
rect 22445 8313 22479 8347
rect 22661 8313 22695 8347
rect 8049 8245 8083 8279
rect 13369 8245 13403 8279
rect 15209 8245 15243 8279
rect 20821 8245 20855 8279
rect 5089 8041 5123 8075
rect 7849 8041 7883 8075
rect 9321 8041 9355 8075
rect 10333 8041 10367 8075
rect 12357 8041 12391 8075
rect 14749 8041 14783 8075
rect 15301 8041 15335 8075
rect 15485 8041 15519 8075
rect 19257 8041 19291 8075
rect 19717 8041 19751 8075
rect 20637 8041 20671 8075
rect 22661 8041 22695 8075
rect 4721 7973 4755 8007
rect 4937 7973 4971 8007
rect 6469 7973 6503 8007
rect 8962 7973 8996 8007
rect 9505 7973 9539 8007
rect 9965 7973 9999 8007
rect 10149 7973 10183 8007
rect 10701 7973 10735 8007
rect 11222 7973 11256 8007
rect 13277 7973 13311 8007
rect 13614 7973 13648 8007
rect 19625 7973 19659 8007
rect 19901 7973 19935 8007
rect 20085 7973 20119 8007
rect 21005 7973 21039 8007
rect 21548 7973 21582 8007
rect 20775 7939 20809 7973
rect 6009 7905 6043 7939
rect 6653 7905 6687 7939
rect 6837 7905 6871 7939
rect 6929 7905 6963 7939
rect 9229 7905 9263 7939
rect 10517 7905 10551 7939
rect 10793 7905 10827 7939
rect 13093 7905 13127 7939
rect 14933 7905 14967 7939
rect 19441 7905 19475 7939
rect 5641 7837 5675 7871
rect 6101 7837 6135 7871
rect 6193 7837 6227 7871
rect 6285 7837 6319 7871
rect 9873 7837 9907 7871
rect 10977 7837 11011 7871
rect 13369 7837 13403 7871
rect 21281 7837 21315 7871
rect 5273 7769 5307 7803
rect 4905 7701 4939 7735
rect 5181 7701 5215 7735
rect 5825 7701 5859 7735
rect 9505 7701 9539 7735
rect 15301 7701 15335 7735
rect 20821 7701 20855 7735
rect 4445 7497 4479 7531
rect 4997 7497 5031 7531
rect 6653 7497 6687 7531
rect 7573 7497 7607 7531
rect 11621 7497 11655 7531
rect 14105 7497 14139 7531
rect 21189 7497 21223 7531
rect 7297 7429 7331 7463
rect 8677 7429 8711 7463
rect 4629 7361 4663 7395
rect 4261 7293 4295 7327
rect 4537 7293 4571 7327
rect 5273 7293 5307 7327
rect 7021 7293 7055 7327
rect 7113 7293 7147 7327
rect 8861 7293 8895 7327
rect 10241 7293 10275 7327
rect 14289 7293 14323 7327
rect 14473 7293 14507 7327
rect 14565 7293 14599 7327
rect 21097 7293 21131 7327
rect 21281 7293 21315 7327
rect 4353 7225 4387 7259
rect 4997 7225 5031 7259
rect 5518 7225 5552 7259
rect 6745 7225 6779 7259
rect 6929 7225 6963 7259
rect 7541 7225 7575 7259
rect 7757 7225 7791 7259
rect 10508 7225 10542 7259
rect 5181 7157 5215 7191
rect 7389 7157 7423 7191
rect 4261 6953 4295 6987
rect 7205 6953 7239 6987
rect 7481 6953 7515 6987
rect 10425 6953 10459 6987
rect 10593 6953 10627 6987
rect 5374 6885 5408 6919
rect 10793 6885 10827 6919
rect 6081 6817 6115 6851
rect 7297 6817 7331 6851
rect 7481 6817 7515 6851
rect 5641 6749 5675 6783
rect 5825 6749 5859 6783
rect 10609 6613 10643 6647
rect 5457 6409 5491 6443
rect 6837 6273 6871 6307
rect 6592 6137 6626 6171
rect 22845 4233 22879 4267
rect 23029 4029 23063 4063
<< metal1 >>
rect 552 23418 23368 23440
rect 552 23366 4322 23418
rect 4374 23366 4386 23418
rect 4438 23366 4450 23418
rect 4502 23366 4514 23418
rect 4566 23366 4578 23418
rect 4630 23366 23368 23418
rect 552 23344 23368 23366
rect 1949 23307 2007 23313
rect 1949 23273 1961 23307
rect 1995 23273 2007 23307
rect 1949 23267 2007 23273
rect 1964 23236 1992 23267
rect 7558 23264 7564 23316
rect 7616 23264 7622 23316
rect 7650 23264 7656 23316
rect 7708 23304 7714 23316
rect 7837 23307 7895 23313
rect 7837 23304 7849 23307
rect 7708 23276 7849 23304
rect 7708 23264 7714 23276
rect 7837 23273 7849 23276
rect 7883 23273 7895 23307
rect 7837 23267 7895 23273
rect 19245 23307 19303 23313
rect 19245 23273 19257 23307
rect 19291 23304 19303 23307
rect 19702 23304 19708 23316
rect 19291 23276 19708 23304
rect 19291 23273 19303 23276
rect 19245 23267 19303 23273
rect 19702 23264 19708 23276
rect 19760 23304 19766 23316
rect 19760 23276 20208 23304
rect 19760 23264 19766 23276
rect 7576 23236 7604 23264
rect 1964 23208 6316 23236
rect 7576 23208 8064 23236
rect 6288 23180 6316 23208
rect 1762 23128 1768 23180
rect 1820 23128 1826 23180
rect 4706 23128 4712 23180
rect 4764 23128 4770 23180
rect 6089 23171 6147 23177
rect 6089 23137 6101 23171
rect 6135 23137 6147 23171
rect 6089 23131 6147 23137
rect 6104 23100 6132 23131
rect 6270 23128 6276 23180
rect 6328 23128 6334 23180
rect 7374 23128 7380 23180
rect 7432 23168 7438 23180
rect 8036 23177 8064 23208
rect 10410 23196 10416 23248
rect 10468 23196 10474 23248
rect 13817 23239 13875 23245
rect 13817 23236 13829 23239
rect 10980 23208 13829 23236
rect 7561 23171 7619 23177
rect 7561 23168 7573 23171
rect 7432 23140 7573 23168
rect 7432 23128 7438 23140
rect 7561 23137 7573 23140
rect 7607 23137 7619 23171
rect 7561 23131 7619 23137
rect 7745 23171 7803 23177
rect 7745 23137 7757 23171
rect 7791 23168 7803 23171
rect 8021 23171 8079 23177
rect 7791 23140 7972 23168
rect 7791 23137 7803 23140
rect 7745 23131 7803 23137
rect 6914 23100 6920 23112
rect 6104 23072 6920 23100
rect 6914 23060 6920 23072
rect 6972 23100 6978 23112
rect 7650 23100 7656 23112
rect 6972 23072 7656 23100
rect 6972 23060 6978 23072
rect 7650 23060 7656 23072
rect 7708 23060 7714 23112
rect 5442 22992 5448 23044
rect 5500 23032 5506 23044
rect 5905 23035 5963 23041
rect 5905 23032 5917 23035
rect 5500 23004 5917 23032
rect 5500 22992 5506 23004
rect 5905 23001 5917 23004
rect 5951 23001 5963 23035
rect 5905 22995 5963 23001
rect 6178 22992 6184 23044
rect 6236 23032 6242 23044
rect 7760 23032 7788 23131
rect 7944 23100 7972 23140
rect 8021 23137 8033 23171
rect 8067 23137 8079 23171
rect 8021 23131 8079 23137
rect 9214 23128 9220 23180
rect 9272 23168 9278 23180
rect 10980 23168 11008 23208
rect 13817 23205 13829 23208
rect 13863 23205 13875 23239
rect 13817 23199 13875 23205
rect 9272 23140 11008 23168
rect 9272 23128 9278 23140
rect 11054 23128 11060 23180
rect 11112 23128 11118 23180
rect 11149 23171 11207 23177
rect 11149 23137 11161 23171
rect 11195 23168 11207 23171
rect 11238 23168 11244 23180
rect 11195 23140 11244 23168
rect 11195 23137 11207 23140
rect 11149 23131 11207 23137
rect 11238 23128 11244 23140
rect 11296 23128 11302 23180
rect 11333 23171 11391 23177
rect 11333 23137 11345 23171
rect 11379 23137 11391 23171
rect 11333 23131 11391 23137
rect 11425 23171 11483 23177
rect 11425 23137 11437 23171
rect 11471 23168 11483 23171
rect 11882 23168 11888 23180
rect 11471 23140 11888 23168
rect 11471 23137 11483 23140
rect 11425 23131 11483 23137
rect 9582 23100 9588 23112
rect 7944 23072 9588 23100
rect 9582 23060 9588 23072
rect 9640 23060 9646 23112
rect 10962 23060 10968 23112
rect 11020 23100 11026 23112
rect 11348 23100 11376 23131
rect 11882 23128 11888 23140
rect 11940 23128 11946 23180
rect 13538 23128 13544 23180
rect 13596 23128 13602 23180
rect 13832 23168 13860 23199
rect 14458 23196 14464 23248
rect 14516 23236 14522 23248
rect 18138 23236 18144 23248
rect 14516 23208 18144 23236
rect 14516 23196 14522 23208
rect 18138 23196 18144 23208
rect 18196 23196 18202 23248
rect 18690 23196 18696 23248
rect 18748 23236 18754 23248
rect 18748 23208 19012 23236
rect 18748 23196 18754 23208
rect 15102 23168 15108 23180
rect 13832 23140 15108 23168
rect 15102 23128 15108 23140
rect 15160 23128 15166 23180
rect 16390 23128 16396 23180
rect 16448 23168 16454 23180
rect 16485 23171 16543 23177
rect 16485 23168 16497 23171
rect 16448 23140 16497 23168
rect 16448 23128 16454 23140
rect 16485 23137 16497 23140
rect 16531 23137 16543 23171
rect 16485 23131 16543 23137
rect 18414 23128 18420 23180
rect 18472 23168 18478 23180
rect 18984 23177 19012 23208
rect 19518 23196 19524 23248
rect 19576 23196 19582 23248
rect 19886 23196 19892 23248
rect 19944 23236 19950 23248
rect 20070 23236 20076 23248
rect 19944 23208 20076 23236
rect 19944 23196 19950 23208
rect 20070 23196 20076 23208
rect 20128 23196 20134 23248
rect 18969 23171 19027 23177
rect 18472 23140 18920 23168
rect 18472 23128 18478 23140
rect 11020 23072 11376 23100
rect 11020 23060 11026 23072
rect 18782 23060 18788 23112
rect 18840 23060 18846 23112
rect 18892 23100 18920 23140
rect 18969 23137 18981 23171
rect 19015 23137 19027 23171
rect 18969 23131 19027 23137
rect 19058 23128 19064 23180
rect 19116 23168 19122 23180
rect 20180 23177 20208 23276
rect 20990 23196 20996 23248
rect 21048 23236 21054 23248
rect 21545 23239 21603 23245
rect 21545 23236 21557 23239
rect 21048 23208 21557 23236
rect 21048 23196 21054 23208
rect 21545 23205 21557 23208
rect 21591 23236 21603 23239
rect 21591 23208 22094 23236
rect 21591 23205 21603 23208
rect 21545 23199 21603 23205
rect 19981 23171 20039 23177
rect 19981 23168 19993 23171
rect 19116 23140 19993 23168
rect 19116 23128 19122 23140
rect 19981 23137 19993 23140
rect 20027 23137 20039 23171
rect 19981 23131 20039 23137
rect 20165 23171 20223 23177
rect 20165 23137 20177 23171
rect 20211 23137 20223 23171
rect 21082 23168 21088 23180
rect 20165 23131 20223 23137
rect 20456 23140 21088 23168
rect 19337 23103 19395 23109
rect 19337 23100 19349 23103
rect 18892 23072 19349 23100
rect 19337 23069 19349 23072
rect 19383 23100 19395 23103
rect 19886 23100 19892 23112
rect 19383 23072 19892 23100
rect 19383 23069 19395 23072
rect 19337 23063 19395 23069
rect 19886 23060 19892 23072
rect 19944 23060 19950 23112
rect 6236 23004 7788 23032
rect 6236 22992 6242 23004
rect 9398 22992 9404 23044
rect 9456 23032 9462 23044
rect 10597 23035 10655 23041
rect 10597 23032 10609 23035
rect 9456 23004 10609 23032
rect 9456 22992 9462 23004
rect 10597 23001 10609 23004
rect 10643 23032 10655 23035
rect 16022 23032 16028 23044
rect 10643 23004 16028 23032
rect 10643 23001 10655 23004
rect 10597 22995 10655 23001
rect 16022 22992 16028 23004
rect 16080 22992 16086 23044
rect 20456 23032 20484 23140
rect 21082 23128 21088 23140
rect 21140 23168 21146 23180
rect 21269 23171 21327 23177
rect 21269 23168 21281 23171
rect 21140 23140 21281 23168
rect 21140 23128 21146 23140
rect 21269 23137 21281 23140
rect 21315 23137 21327 23171
rect 21269 23131 21327 23137
rect 21358 23128 21364 23180
rect 21416 23128 21422 23180
rect 21450 23128 21456 23180
rect 21508 23168 21514 23180
rect 21637 23171 21695 23177
rect 21637 23168 21649 23171
rect 21508 23140 21649 23168
rect 21508 23128 21514 23140
rect 21637 23137 21649 23140
rect 21683 23137 21695 23171
rect 21637 23131 21695 23137
rect 21729 23171 21787 23177
rect 21729 23137 21741 23171
rect 21775 23137 21787 23171
rect 21729 23131 21787 23137
rect 20530 23060 20536 23112
rect 20588 23100 20594 23112
rect 21744 23100 21772 23131
rect 21910 23128 21916 23180
rect 21968 23128 21974 23180
rect 20588 23072 21772 23100
rect 20588 23060 20594 23072
rect 17512 23004 20484 23032
rect 22066 23032 22094 23208
rect 22278 23128 22284 23180
rect 22336 23168 22342 23180
rect 22373 23171 22431 23177
rect 22373 23168 22385 23171
rect 22336 23140 22385 23168
rect 22336 23128 22342 23140
rect 22373 23137 22385 23140
rect 22419 23137 22431 23171
rect 22373 23131 22431 23137
rect 22557 23103 22615 23109
rect 22557 23069 22569 23103
rect 22603 23069 22615 23103
rect 22557 23063 22615 23069
rect 22572 23032 22600 23063
rect 22066 23004 22600 23032
rect 17512 22976 17540 23004
rect 4890 22924 4896 22976
rect 4948 22924 4954 22976
rect 5350 22924 5356 22976
rect 5408 22964 5414 22976
rect 6457 22967 6515 22973
rect 6457 22964 6469 22967
rect 5408 22936 6469 22964
rect 5408 22924 5414 22936
rect 6457 22933 6469 22936
rect 6503 22933 6515 22967
rect 6457 22927 6515 22933
rect 7653 22967 7711 22973
rect 7653 22933 7665 22967
rect 7699 22964 7711 22967
rect 7742 22964 7748 22976
rect 7699 22936 7748 22964
rect 7699 22933 7711 22936
rect 7653 22927 7711 22933
rect 7742 22924 7748 22936
rect 7800 22924 7806 22976
rect 11609 22967 11667 22973
rect 11609 22933 11621 22967
rect 11655 22964 11667 22967
rect 13538 22964 13544 22976
rect 11655 22936 13544 22964
rect 11655 22933 11667 22936
rect 11609 22927 11667 22933
rect 13538 22924 13544 22936
rect 13596 22964 13602 22976
rect 14274 22964 14280 22976
rect 13596 22936 14280 22964
rect 13596 22924 13602 22936
rect 14274 22924 14280 22936
rect 14332 22924 14338 22976
rect 16669 22967 16727 22973
rect 16669 22933 16681 22967
rect 16715 22964 16727 22967
rect 17494 22964 17500 22976
rect 16715 22936 17500 22964
rect 16715 22933 16727 22936
rect 16669 22927 16727 22933
rect 17494 22924 17500 22936
rect 17552 22924 17558 22976
rect 19978 22924 19984 22976
rect 20036 22924 20042 22976
rect 20070 22924 20076 22976
rect 20128 22964 20134 22976
rect 21358 22964 21364 22976
rect 20128 22936 21364 22964
rect 20128 22924 20134 22936
rect 21358 22924 21364 22936
rect 21416 22924 21422 22976
rect 21453 22967 21511 22973
rect 21453 22933 21465 22967
rect 21499 22964 21511 22967
rect 21726 22964 21732 22976
rect 21499 22936 21732 22964
rect 21499 22933 21511 22936
rect 21453 22927 21511 22933
rect 21726 22924 21732 22936
rect 21784 22924 21790 22976
rect 21913 22967 21971 22973
rect 21913 22933 21925 22967
rect 21959 22964 21971 22967
rect 22554 22964 22560 22976
rect 21959 22936 22560 22964
rect 21959 22933 21971 22936
rect 21913 22927 21971 22933
rect 22554 22924 22560 22936
rect 22612 22924 22618 22976
rect 552 22874 23368 22896
rect 552 22822 3662 22874
rect 3714 22822 3726 22874
rect 3778 22822 3790 22874
rect 3842 22822 3854 22874
rect 3906 22822 3918 22874
rect 3970 22822 23368 22874
rect 552 22800 23368 22822
rect 5077 22763 5135 22769
rect 5077 22729 5089 22763
rect 5123 22729 5135 22763
rect 5077 22723 5135 22729
rect 5092 22692 5120 22723
rect 9766 22720 9772 22772
rect 9824 22760 9830 22772
rect 9861 22763 9919 22769
rect 9861 22760 9873 22763
rect 9824 22732 9873 22760
rect 9824 22720 9830 22732
rect 9861 22729 9873 22732
rect 9907 22729 9919 22763
rect 10410 22760 10416 22772
rect 9861 22723 9919 22729
rect 9968 22732 10416 22760
rect 9968 22704 9996 22732
rect 10410 22720 10416 22732
rect 10468 22720 10474 22772
rect 13173 22763 13231 22769
rect 13173 22729 13185 22763
rect 13219 22760 13231 22763
rect 13998 22760 14004 22772
rect 13219 22732 14004 22760
rect 13219 22729 13231 22732
rect 13173 22723 13231 22729
rect 13998 22720 14004 22732
rect 14056 22720 14062 22772
rect 14274 22720 14280 22772
rect 14332 22720 14338 22772
rect 15194 22720 15200 22772
rect 15252 22760 15258 22772
rect 15289 22763 15347 22769
rect 15289 22760 15301 22763
rect 15252 22732 15301 22760
rect 15252 22720 15258 22732
rect 15289 22729 15301 22732
rect 15335 22760 15347 22763
rect 16390 22760 16396 22772
rect 15335 22732 16396 22760
rect 15335 22729 15347 22732
rect 15289 22723 15347 22729
rect 5350 22692 5356 22704
rect 5092 22664 5356 22692
rect 5350 22652 5356 22664
rect 5408 22692 5414 22704
rect 5537 22695 5595 22701
rect 5537 22692 5549 22695
rect 5408 22664 5549 22692
rect 5408 22652 5414 22664
rect 5537 22661 5549 22664
rect 5583 22661 5595 22695
rect 5537 22655 5595 22661
rect 7374 22652 7380 22704
rect 7432 22692 7438 22704
rect 9950 22692 9956 22704
rect 7432 22664 9956 22692
rect 7432 22652 7438 22664
rect 9950 22652 9956 22664
rect 10008 22652 10014 22704
rect 10137 22695 10195 22701
rect 10137 22661 10149 22695
rect 10183 22692 10195 22695
rect 11054 22692 11060 22704
rect 10183 22664 11060 22692
rect 10183 22661 10195 22664
rect 10137 22655 10195 22661
rect 11054 22652 11060 22664
rect 11112 22652 11118 22704
rect 12805 22695 12863 22701
rect 12805 22661 12817 22695
rect 12851 22661 12863 22695
rect 13906 22692 13912 22704
rect 12805 22655 12863 22661
rect 13372 22664 13912 22692
rect 4890 22584 4896 22636
rect 4948 22624 4954 22636
rect 5626 22624 5632 22636
rect 4948 22596 5632 22624
rect 4948 22584 4954 22596
rect 5626 22584 5632 22596
rect 5684 22624 5690 22636
rect 5684 22596 5764 22624
rect 5684 22584 5690 22596
rect 5353 22559 5411 22565
rect 5353 22525 5365 22559
rect 5399 22525 5411 22559
rect 5353 22519 5411 22525
rect 4890 22448 4896 22500
rect 4948 22448 4954 22500
rect 5368 22488 5396 22519
rect 5442 22516 5448 22568
rect 5500 22516 5506 22568
rect 5736 22565 5764 22596
rect 9398 22584 9404 22636
rect 9456 22584 9462 22636
rect 10962 22624 10968 22636
rect 9692 22596 10364 22624
rect 5721 22559 5779 22565
rect 5721 22525 5733 22559
rect 5767 22525 5779 22559
rect 5721 22519 5779 22525
rect 6362 22516 6368 22568
rect 6420 22516 6426 22568
rect 7190 22516 7196 22568
rect 7248 22556 7254 22568
rect 8389 22559 8447 22565
rect 8389 22556 8401 22559
rect 7248 22528 8401 22556
rect 7248 22516 7254 22528
rect 8389 22525 8401 22528
rect 8435 22556 8447 22559
rect 9214 22556 9220 22568
rect 8435 22528 9220 22556
rect 8435 22525 8447 22528
rect 8389 22519 8447 22525
rect 9214 22516 9220 22528
rect 9272 22516 9278 22568
rect 5994 22488 6000 22500
rect 5368 22460 6000 22488
rect 5994 22448 6000 22460
rect 6052 22448 6058 22500
rect 6178 22448 6184 22500
rect 6236 22448 6242 22500
rect 7650 22448 7656 22500
rect 7708 22448 7714 22500
rect 9582 22448 9588 22500
rect 9640 22488 9646 22500
rect 9692 22497 9720 22596
rect 9677 22491 9735 22497
rect 9677 22488 9689 22491
rect 9640 22460 9689 22488
rect 9640 22448 9646 22460
rect 9677 22457 9689 22460
rect 9723 22457 9735 22491
rect 9677 22451 9735 22457
rect 9766 22448 9772 22500
rect 9824 22488 9830 22500
rect 10336 22497 10364 22596
rect 10428 22596 10968 22624
rect 10428 22568 10456 22596
rect 10962 22584 10968 22596
rect 11020 22624 11026 22636
rect 11333 22627 11391 22633
rect 11333 22624 11345 22627
rect 11020 22596 11345 22624
rect 11020 22584 11026 22596
rect 11333 22593 11345 22596
rect 11379 22593 11391 22627
rect 11333 22587 11391 22593
rect 11517 22627 11575 22633
rect 11517 22593 11529 22627
rect 11563 22624 11575 22627
rect 12820 22624 12848 22655
rect 13081 22627 13139 22633
rect 13081 22624 13093 22627
rect 11563 22596 12020 22624
rect 12820 22596 13093 22624
rect 11563 22593 11575 22596
rect 11517 22587 11575 22593
rect 10410 22516 10416 22568
rect 10468 22516 10474 22568
rect 11241 22559 11299 22565
rect 11241 22525 11253 22559
rect 11287 22525 11299 22559
rect 11241 22519 11299 22525
rect 10137 22491 10195 22497
rect 10137 22488 10149 22491
rect 9824 22460 10149 22488
rect 9824 22448 9830 22460
rect 10137 22457 10149 22460
rect 10183 22457 10195 22491
rect 10137 22451 10195 22457
rect 10321 22491 10379 22497
rect 10321 22457 10333 22491
rect 10367 22488 10379 22491
rect 11054 22488 11060 22500
rect 10367 22460 11060 22488
rect 10367 22457 10379 22460
rect 10321 22451 10379 22457
rect 11054 22448 11060 22460
rect 11112 22488 11118 22500
rect 11256 22488 11284 22519
rect 11606 22516 11612 22568
rect 11664 22516 11670 22568
rect 11701 22559 11759 22565
rect 11701 22525 11713 22559
rect 11747 22525 11759 22559
rect 11701 22519 11759 22525
rect 11112 22460 11284 22488
rect 11112 22448 11118 22460
rect 11514 22448 11520 22500
rect 11572 22488 11578 22500
rect 11716 22488 11744 22519
rect 11882 22516 11888 22568
rect 11940 22516 11946 22568
rect 11992 22565 12020 22596
rect 13081 22593 13093 22596
rect 13127 22624 13139 22627
rect 13170 22624 13176 22636
rect 13127 22596 13176 22624
rect 13127 22593 13139 22596
rect 13081 22587 13139 22593
rect 13170 22584 13176 22596
rect 13228 22584 13234 22636
rect 11977 22559 12035 22565
rect 11977 22525 11989 22559
rect 12023 22556 12035 22559
rect 12066 22556 12072 22568
rect 12023 22528 12072 22556
rect 12023 22525 12035 22528
rect 11977 22519 12035 22525
rect 12066 22516 12072 22528
rect 12124 22516 12130 22568
rect 12161 22559 12219 22565
rect 12161 22525 12173 22559
rect 12207 22556 12219 22559
rect 12250 22556 12256 22568
rect 12207 22528 12256 22556
rect 12207 22525 12219 22528
rect 12161 22519 12219 22525
rect 12250 22516 12256 22528
rect 12308 22556 12314 22568
rect 12529 22559 12587 22565
rect 12529 22556 12541 22559
rect 12308 22528 12541 22556
rect 12308 22516 12314 22528
rect 12529 22525 12541 22528
rect 12575 22525 12587 22559
rect 12529 22519 12587 22525
rect 12621 22559 12679 22565
rect 12621 22525 12633 22559
rect 12667 22556 12679 22559
rect 12667 22528 13216 22556
rect 12667 22525 12679 22528
rect 12621 22519 12679 22525
rect 11572 22460 11744 22488
rect 11572 22448 11578 22460
rect 12802 22448 12808 22500
rect 12860 22448 12866 22500
rect 13188 22488 13216 22528
rect 13262 22516 13268 22568
rect 13320 22516 13326 22568
rect 13372 22565 13400 22664
rect 13906 22652 13912 22664
rect 13964 22692 13970 22704
rect 14093 22695 14151 22701
rect 14093 22692 14105 22695
rect 13964 22664 14105 22692
rect 13964 22652 13970 22664
rect 14093 22661 14105 22664
rect 14139 22661 14151 22695
rect 14093 22655 14151 22661
rect 15473 22695 15531 22701
rect 15473 22661 15485 22695
rect 15519 22692 15531 22695
rect 15746 22692 15752 22704
rect 15519 22664 15752 22692
rect 15519 22661 15531 22664
rect 15473 22655 15531 22661
rect 15746 22652 15752 22664
rect 15804 22652 15810 22704
rect 13538 22584 13544 22636
rect 13596 22584 13602 22636
rect 13725 22627 13783 22633
rect 13725 22593 13737 22627
rect 13771 22624 13783 22627
rect 13814 22624 13820 22636
rect 13771 22596 13820 22624
rect 13771 22593 13783 22596
rect 13725 22587 13783 22593
rect 13814 22584 13820 22596
rect 13872 22624 13878 22636
rect 15856 22633 15884 22732
rect 16390 22720 16396 22732
rect 16448 22720 16454 22772
rect 18325 22763 18383 22769
rect 18325 22729 18337 22763
rect 18371 22729 18383 22763
rect 18325 22723 18383 22729
rect 18509 22763 18567 22769
rect 18509 22729 18521 22763
rect 18555 22760 18567 22763
rect 19058 22760 19064 22772
rect 18555 22732 19064 22760
rect 18555 22729 18567 22732
rect 18509 22723 18567 22729
rect 16485 22695 16543 22701
rect 16485 22661 16497 22695
rect 16531 22692 16543 22695
rect 16758 22692 16764 22704
rect 16531 22664 16764 22692
rect 16531 22661 16543 22664
rect 16485 22655 16543 22661
rect 16758 22652 16764 22664
rect 16816 22652 16822 22704
rect 16850 22652 16856 22704
rect 16908 22692 16914 22704
rect 18340 22692 18368 22723
rect 19058 22720 19064 22732
rect 19116 22720 19122 22772
rect 20717 22763 20775 22769
rect 20717 22729 20729 22763
rect 20763 22760 20775 22763
rect 21450 22760 21456 22772
rect 20763 22732 21456 22760
rect 20763 22729 20775 22732
rect 20717 22723 20775 22729
rect 18782 22692 18788 22704
rect 16908 22664 18788 22692
rect 16908 22652 16914 22664
rect 18782 22652 18788 22664
rect 18840 22652 18846 22704
rect 20732 22692 20760 22723
rect 21450 22720 21456 22732
rect 21508 22720 21514 22772
rect 21545 22763 21603 22769
rect 21545 22729 21557 22763
rect 21591 22760 21603 22763
rect 21910 22760 21916 22772
rect 21591 22732 21916 22760
rect 21591 22729 21603 22732
rect 21545 22723 21603 22729
rect 19260 22664 20760 22692
rect 15841 22627 15899 22633
rect 13872 22596 14596 22624
rect 13872 22584 13878 22596
rect 13357 22559 13415 22565
rect 13357 22525 13369 22559
rect 13403 22525 13415 22559
rect 13357 22519 13415 22525
rect 13630 22516 13636 22568
rect 13688 22556 13694 22568
rect 14568 22565 14596 22596
rect 15841 22593 15853 22627
rect 15887 22593 15899 22627
rect 15841 22587 15899 22593
rect 16022 22584 16028 22636
rect 16080 22624 16086 22636
rect 18690 22624 18696 22636
rect 16080 22596 18696 22624
rect 16080 22584 16086 22596
rect 14001 22559 14059 22565
rect 14001 22556 14013 22559
rect 13688 22528 14013 22556
rect 13688 22516 13694 22528
rect 14001 22525 14013 22528
rect 14047 22556 14059 22559
rect 14553 22559 14611 22565
rect 14047 22528 14290 22556
rect 14047 22525 14059 22528
rect 14001 22519 14059 22525
rect 14231 22525 14290 22528
rect 13446 22488 13452 22500
rect 13188 22460 13452 22488
rect 13446 22448 13452 22460
rect 13504 22448 13510 22500
rect 14231 22491 14243 22525
rect 14277 22494 14290 22525
rect 14553 22525 14565 22559
rect 14599 22525 14611 22559
rect 14553 22519 14611 22525
rect 14642 22516 14648 22568
rect 14700 22556 14706 22568
rect 15933 22559 15991 22565
rect 14700 22528 14745 22556
rect 15120 22528 15608 22556
rect 14700 22516 14706 22528
rect 15120 22500 15148 22528
rect 14277 22491 14289 22494
rect 14231 22485 14289 22491
rect 14458 22448 14464 22500
rect 14516 22448 14522 22500
rect 15102 22448 15108 22500
rect 15160 22448 15166 22500
rect 15580 22488 15608 22528
rect 15933 22525 15945 22559
rect 15979 22552 15991 22559
rect 16040 22552 16068 22584
rect 15979 22525 16068 22552
rect 15933 22524 16068 22525
rect 16209 22559 16267 22565
rect 16209 22525 16221 22559
rect 16255 22556 16267 22559
rect 16390 22556 16396 22568
rect 16255 22528 16396 22556
rect 16255 22525 16267 22528
rect 15933 22519 15991 22524
rect 16209 22519 16267 22525
rect 16390 22516 16396 22528
rect 16448 22516 16454 22568
rect 16500 22528 17908 22556
rect 16500 22500 16528 22528
rect 15580 22460 16344 22488
rect 5074 22380 5080 22432
rect 5132 22420 5138 22432
rect 5442 22420 5448 22432
rect 5132 22392 5448 22420
rect 5132 22380 5138 22392
rect 5442 22380 5448 22392
rect 5500 22380 5506 22432
rect 8478 22380 8484 22432
rect 8536 22380 8542 22432
rect 9030 22380 9036 22432
rect 9088 22380 9094 22432
rect 9858 22380 9864 22432
rect 9916 22429 9922 22432
rect 9916 22423 9935 22429
rect 9923 22389 9935 22423
rect 9916 22383 9935 22389
rect 9916 22380 9922 22383
rect 10042 22380 10048 22432
rect 10100 22380 10106 22432
rect 10873 22423 10931 22429
rect 10873 22389 10885 22423
rect 10919 22420 10931 22423
rect 11422 22420 11428 22432
rect 10919 22392 11428 22420
rect 10919 22389 10931 22392
rect 10873 22383 10931 22389
rect 11422 22380 11428 22392
rect 11480 22380 11486 22432
rect 13354 22380 13360 22432
rect 13412 22420 13418 22432
rect 13909 22423 13967 22429
rect 13909 22420 13921 22423
rect 13412 22392 13921 22420
rect 13412 22380 13418 22392
rect 13909 22389 13921 22392
rect 13955 22420 13967 22423
rect 14476 22420 14504 22448
rect 16316 22432 16344 22460
rect 16482 22448 16488 22500
rect 16540 22448 16546 22500
rect 16761 22491 16819 22497
rect 16761 22457 16773 22491
rect 16807 22488 16819 22491
rect 16850 22488 16856 22500
rect 16807 22460 16856 22488
rect 16807 22457 16819 22460
rect 16761 22451 16819 22457
rect 13955 22392 14504 22420
rect 13955 22389 13967 22392
rect 13909 22383 13967 22389
rect 14918 22380 14924 22432
rect 14976 22380 14982 22432
rect 15286 22380 15292 22432
rect 15344 22429 15350 22432
rect 15344 22423 15363 22429
rect 15351 22389 15363 22423
rect 15344 22383 15363 22389
rect 15565 22423 15623 22429
rect 15565 22389 15577 22423
rect 15611 22420 15623 22423
rect 15746 22420 15752 22432
rect 15611 22392 15752 22420
rect 15611 22389 15623 22392
rect 15565 22383 15623 22389
rect 15344 22380 15350 22383
rect 15746 22380 15752 22392
rect 15804 22380 15810 22432
rect 16298 22380 16304 22432
rect 16356 22380 16362 22432
rect 16390 22380 16396 22432
rect 16448 22420 16454 22432
rect 16776 22420 16804 22451
rect 16850 22448 16856 22460
rect 16908 22448 16914 22500
rect 17494 22448 17500 22500
rect 17552 22448 17558 22500
rect 17586 22448 17592 22500
rect 17644 22448 17650 22500
rect 17770 22448 17776 22500
rect 17828 22448 17834 22500
rect 17880 22488 17908 22528
rect 18156 22497 18184 22596
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 18800 22556 18828 22652
rect 19260 22636 19288 22664
rect 19242 22584 19248 22636
rect 19300 22584 19306 22636
rect 19352 22596 19932 22624
rect 19352 22556 19380 22596
rect 18371 22525 18429 22531
rect 18800 22528 19380 22556
rect 18371 22522 18383 22525
rect 18141 22491 18199 22497
rect 17880 22460 18092 22488
rect 16448 22392 16804 22420
rect 16448 22380 16454 22392
rect 17954 22380 17960 22432
rect 18012 22380 18018 22432
rect 18064 22420 18092 22460
rect 18141 22457 18153 22491
rect 18187 22457 18199 22491
rect 18356 22491 18383 22522
rect 18417 22500 18429 22525
rect 19794 22516 19800 22568
rect 19852 22516 19858 22568
rect 19904 22556 19932 22596
rect 19978 22584 19984 22636
rect 20036 22584 20042 22636
rect 20990 22584 20996 22636
rect 21048 22624 21054 22636
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 21048 22596 21097 22624
rect 21048 22584 21054 22596
rect 21085 22593 21097 22596
rect 21131 22593 21143 22627
rect 21085 22587 21143 22593
rect 21177 22559 21235 22565
rect 21177 22556 21189 22559
rect 19904 22528 21189 22556
rect 21177 22525 21189 22528
rect 21223 22525 21235 22559
rect 21177 22519 21235 22525
rect 18417 22491 18420 22500
rect 18356 22488 18420 22491
rect 18141 22451 18199 22457
rect 18248 22460 18420 22488
rect 18248 22420 18276 22460
rect 18414 22448 18420 22460
rect 18472 22448 18478 22500
rect 18693 22491 18751 22497
rect 18693 22457 18705 22491
rect 18739 22488 18751 22491
rect 18782 22488 18788 22500
rect 18739 22460 18788 22488
rect 18739 22457 18751 22460
rect 18693 22451 18751 22457
rect 18782 22448 18788 22460
rect 18840 22448 18846 22500
rect 18874 22448 18880 22500
rect 18932 22448 18938 22500
rect 18966 22448 18972 22500
rect 19024 22488 19030 22500
rect 20530 22488 20536 22500
rect 19024 22460 20536 22488
rect 19024 22448 19030 22460
rect 20530 22448 20536 22460
rect 20588 22448 20594 22500
rect 20749 22491 20807 22497
rect 20749 22457 20761 22491
rect 20795 22488 20807 22491
rect 21560 22488 21588 22723
rect 21910 22720 21916 22732
rect 21968 22720 21974 22772
rect 21821 22695 21879 22701
rect 21821 22661 21833 22695
rect 21867 22692 21879 22695
rect 22002 22692 22008 22704
rect 21867 22664 22008 22692
rect 21867 22661 21879 22664
rect 21821 22655 21879 22661
rect 22002 22652 22008 22664
rect 22060 22652 22066 22704
rect 20795 22460 21588 22488
rect 22097 22491 22155 22497
rect 20795 22457 20807 22460
rect 20749 22451 20807 22457
rect 22097 22457 22109 22491
rect 22143 22488 22155 22491
rect 22186 22488 22192 22500
rect 22143 22460 22192 22488
rect 22143 22457 22155 22460
rect 22097 22451 22155 22457
rect 22186 22448 22192 22460
rect 22244 22448 22250 22500
rect 18064 22392 18276 22420
rect 19058 22380 19064 22432
rect 19116 22380 19122 22432
rect 20901 22423 20959 22429
rect 20901 22389 20913 22423
rect 20947 22420 20959 22423
rect 21542 22420 21548 22432
rect 20947 22392 21548 22420
rect 20947 22389 20959 22392
rect 20901 22383 20959 22389
rect 21542 22380 21548 22392
rect 21600 22380 21606 22432
rect 21634 22380 21640 22432
rect 21692 22380 21698 22432
rect 552 22330 23368 22352
rect 552 22278 4322 22330
rect 4374 22278 4386 22330
rect 4438 22278 4450 22330
rect 4502 22278 4514 22330
rect 4566 22278 4578 22330
rect 4630 22278 23368 22330
rect 552 22256 23368 22278
rect 11606 22176 11612 22228
rect 11664 22216 11670 22228
rect 12713 22219 12771 22225
rect 11664 22188 12388 22216
rect 11664 22176 11670 22188
rect 7558 22108 7564 22160
rect 7616 22148 7622 22160
rect 9214 22148 9220 22160
rect 7616 22120 7788 22148
rect 7616 22108 7622 22120
rect 5445 22083 5503 22089
rect 5445 22049 5457 22083
rect 5491 22080 5503 22083
rect 5626 22080 5632 22092
rect 5491 22052 5632 22080
rect 5491 22049 5503 22052
rect 5445 22043 5503 22049
rect 5626 22040 5632 22052
rect 5684 22080 5690 22092
rect 5905 22083 5963 22089
rect 5905 22080 5917 22083
rect 5684 22052 5917 22080
rect 5684 22040 5690 22052
rect 5905 22049 5917 22052
rect 5951 22049 5963 22083
rect 5905 22043 5963 22049
rect 6270 22040 6276 22092
rect 6328 22040 6334 22092
rect 6549 22083 6607 22089
rect 6549 22049 6561 22083
rect 6595 22080 6607 22083
rect 6914 22080 6920 22092
rect 6595 22052 6920 22080
rect 6595 22049 6607 22052
rect 6549 22043 6607 22049
rect 6914 22040 6920 22052
rect 6972 22040 6978 22092
rect 7760 22089 7788 22120
rect 8956 22120 9220 22148
rect 8956 22114 8984 22120
rect 7745 22083 7803 22089
rect 7745 22080 7757 22083
rect 7723 22052 7757 22080
rect 7745 22049 7757 22052
rect 7791 22049 7803 22083
rect 7745 22043 7803 22049
rect 8202 22040 8208 22092
rect 8260 22080 8266 22092
rect 8864 22089 8984 22114
rect 9214 22108 9220 22120
rect 9272 22108 9278 22160
rect 10042 22108 10048 22160
rect 10100 22148 10106 22160
rect 10689 22151 10747 22157
rect 10689 22148 10701 22151
rect 10100 22120 10701 22148
rect 10100 22108 10106 22120
rect 10689 22117 10701 22120
rect 10735 22148 10747 22151
rect 11238 22148 11244 22160
rect 10735 22120 11244 22148
rect 10735 22117 10747 22120
rect 10689 22111 10747 22117
rect 11238 22108 11244 22120
rect 11296 22148 11302 22160
rect 11882 22148 11888 22160
rect 11296 22120 11468 22148
rect 11296 22108 11302 22120
rect 8481 22083 8539 22089
rect 8481 22080 8493 22083
rect 8260 22052 8493 22080
rect 8260 22040 8266 22052
rect 8481 22049 8493 22052
rect 8527 22049 8539 22083
rect 8849 22086 8984 22089
rect 8849 22083 8907 22086
rect 8849 22080 8861 22083
rect 8827 22052 8861 22080
rect 8481 22043 8539 22049
rect 8849 22049 8861 22052
rect 8895 22049 8907 22083
rect 8849 22043 8907 22049
rect 9033 22083 9091 22089
rect 9033 22049 9045 22083
rect 9079 22049 9091 22083
rect 9033 22043 9091 22049
rect 9585 22083 9643 22089
rect 9585 22049 9597 22083
rect 9631 22080 9643 22083
rect 9858 22080 9864 22092
rect 9631 22052 9864 22080
rect 9631 22049 9643 22052
rect 9585 22043 9643 22049
rect 9048 22012 9076 22043
rect 9858 22040 9864 22052
rect 9916 22080 9922 22092
rect 10321 22083 10379 22089
rect 10321 22080 10333 22083
rect 9916 22052 10333 22080
rect 9916 22040 9922 22052
rect 10321 22049 10333 22052
rect 10367 22049 10379 22083
rect 10321 22043 10379 22049
rect 10505 22083 10563 22089
rect 10505 22049 10517 22083
rect 10551 22049 10563 22083
rect 10505 22043 10563 22049
rect 8864 21984 9076 22012
rect 5997 21947 6055 21953
rect 5997 21913 6009 21947
rect 6043 21944 6055 21947
rect 7374 21944 7380 21956
rect 6043 21916 7380 21944
rect 6043 21913 6055 21916
rect 5997 21907 6055 21913
rect 7374 21904 7380 21916
rect 7432 21904 7438 21956
rect 7466 21904 7472 21956
rect 7524 21904 7530 21956
rect 7650 21904 7656 21956
rect 7708 21944 7714 21956
rect 8202 21944 8208 21956
rect 7708 21916 8208 21944
rect 7708 21904 7714 21916
rect 8202 21904 8208 21916
rect 8260 21904 8266 21956
rect 5258 21836 5264 21888
rect 5316 21836 5322 21888
rect 6362 21836 6368 21888
rect 6420 21876 6426 21888
rect 8864 21876 8892 21984
rect 9214 21972 9220 22024
rect 9272 22012 9278 22024
rect 9309 22015 9367 22021
rect 9309 22012 9321 22015
rect 9272 21984 9321 22012
rect 9272 21972 9278 21984
rect 9309 21981 9321 21984
rect 9355 21981 9367 22015
rect 9309 21975 9367 21981
rect 10226 21972 10232 22024
rect 10284 21972 10290 22024
rect 8941 21947 8999 21953
rect 8941 21913 8953 21947
rect 8987 21944 8999 21947
rect 9674 21944 9680 21956
rect 8987 21916 9680 21944
rect 8987 21913 8999 21916
rect 8941 21907 8999 21913
rect 9674 21904 9680 21916
rect 9732 21904 9738 21956
rect 10134 21904 10140 21956
rect 10192 21944 10198 21956
rect 10520 21944 10548 22043
rect 11146 22040 11152 22092
rect 11204 22040 11210 22092
rect 11440 22089 11468 22120
rect 11716 22120 11888 22148
rect 11425 22083 11483 22089
rect 11425 22049 11437 22083
rect 11471 22049 11483 22083
rect 11716 22080 11744 22120
rect 11882 22108 11888 22120
rect 11940 22148 11946 22160
rect 11940 22120 12296 22148
rect 11940 22108 11946 22120
rect 11790 22080 11796 22092
rect 11716 22052 11796 22080
rect 11425 22043 11483 22049
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 12066 22040 12072 22092
rect 12124 22040 12130 22092
rect 12268 22089 12296 22120
rect 12360 22089 12388 22188
rect 12713 22185 12725 22219
rect 12759 22216 12771 22219
rect 12802 22216 12808 22228
rect 12759 22188 12808 22216
rect 12759 22185 12771 22188
rect 12713 22179 12771 22185
rect 12802 22176 12808 22188
rect 12860 22176 12866 22228
rect 14918 22176 14924 22228
rect 14976 22216 14982 22228
rect 15473 22219 15531 22225
rect 15473 22216 15485 22219
rect 14976 22188 15485 22216
rect 14976 22176 14982 22188
rect 15473 22185 15485 22188
rect 15519 22185 15531 22219
rect 15473 22179 15531 22185
rect 16298 22176 16304 22228
rect 16356 22216 16362 22228
rect 16356 22188 17816 22216
rect 16356 22176 16362 22188
rect 13096 22120 13584 22148
rect 12253 22083 12311 22089
rect 12253 22080 12265 22083
rect 12231 22052 12265 22080
rect 12253 22049 12265 22052
rect 12299 22049 12311 22083
rect 12253 22043 12311 22049
rect 12345 22083 12403 22089
rect 12345 22049 12357 22083
rect 12391 22049 12403 22083
rect 12345 22043 12403 22049
rect 12437 22083 12495 22089
rect 12437 22049 12449 22083
rect 12483 22049 12495 22083
rect 12437 22043 12495 22049
rect 10962 21972 10968 22024
rect 11020 22012 11026 22024
rect 11977 22015 12035 22021
rect 11977 22012 11989 22015
rect 11020 21984 11989 22012
rect 11020 21972 11026 21984
rect 11977 21981 11989 21984
rect 12023 21981 12035 22015
rect 12452 22012 12480 22043
rect 12710 22040 12716 22092
rect 12768 22080 12774 22092
rect 13096 22080 13124 22120
rect 12768 22052 13124 22080
rect 13173 22083 13231 22089
rect 12768 22040 12774 22052
rect 13173 22049 13185 22083
rect 13219 22080 13231 22083
rect 13446 22080 13452 22092
rect 13219 22052 13452 22080
rect 13219 22049 13231 22052
rect 13173 22043 13231 22049
rect 13446 22040 13452 22052
rect 13504 22040 13510 22092
rect 13556 22080 13584 22120
rect 15562 22108 15568 22160
rect 15620 22108 15626 22160
rect 15933 22151 15991 22157
rect 15933 22117 15945 22151
rect 15979 22148 15991 22151
rect 17034 22148 17040 22160
rect 15979 22120 17040 22148
rect 15979 22117 15991 22120
rect 15933 22111 15991 22117
rect 17034 22108 17040 22120
rect 17092 22148 17098 22160
rect 17092 22120 17632 22148
rect 17092 22108 17098 22120
rect 13556 22052 14044 22080
rect 11977 21975 12035 21981
rect 12084 21984 12480 22012
rect 11330 21944 11336 21956
rect 10192 21916 11336 21944
rect 10192 21904 10198 21916
rect 11330 21904 11336 21916
rect 11388 21944 11394 21956
rect 12084 21944 12112 21984
rect 13078 21972 13084 22024
rect 13136 21972 13142 22024
rect 13814 21972 13820 22024
rect 13872 21972 13878 22024
rect 14016 22012 14044 22052
rect 14090 22040 14096 22092
rect 14148 22080 14154 22092
rect 14642 22080 14648 22092
rect 14148 22052 14648 22080
rect 14148 22040 14154 22052
rect 14642 22040 14648 22052
rect 14700 22040 14706 22092
rect 15746 22040 15752 22092
rect 15804 22040 15810 22092
rect 16114 22040 16120 22092
rect 16172 22040 16178 22092
rect 16574 22040 16580 22092
rect 16632 22040 16638 22092
rect 16758 22040 16764 22092
rect 16816 22080 16822 22092
rect 16945 22083 17003 22089
rect 16945 22080 16957 22083
rect 16816 22052 16957 22080
rect 16816 22040 16822 22052
rect 16945 22049 16957 22052
rect 16991 22080 17003 22083
rect 17126 22080 17132 22092
rect 16991 22052 17132 22080
rect 16991 22049 17003 22052
rect 16945 22043 17003 22049
rect 17126 22040 17132 22052
rect 17184 22040 17190 22092
rect 17402 22040 17408 22092
rect 17460 22040 17466 22092
rect 17497 22083 17555 22089
rect 17497 22049 17509 22083
rect 17543 22049 17555 22083
rect 17604 22080 17632 22120
rect 17674 22083 17732 22089
rect 17674 22080 17686 22083
rect 17604 22052 17686 22080
rect 17497 22043 17555 22049
rect 17674 22049 17686 22052
rect 17720 22049 17732 22083
rect 17788 22080 17816 22188
rect 18230 22176 18236 22228
rect 18288 22216 18294 22228
rect 18325 22219 18383 22225
rect 18325 22216 18337 22219
rect 18288 22188 18337 22216
rect 18288 22176 18294 22188
rect 18325 22185 18337 22188
rect 18371 22216 18383 22219
rect 18617 22219 18675 22225
rect 18617 22216 18629 22219
rect 18371 22188 18629 22216
rect 18371 22185 18383 22188
rect 18325 22179 18383 22185
rect 18617 22185 18629 22188
rect 18663 22185 18675 22219
rect 18617 22179 18675 22185
rect 18782 22176 18788 22228
rect 18840 22176 18846 22228
rect 21542 22176 21548 22228
rect 21600 22216 21606 22228
rect 21600 22188 22324 22216
rect 21600 22176 21606 22188
rect 18414 22108 18420 22160
rect 18472 22108 18478 22160
rect 21269 22151 21327 22157
rect 21269 22117 21281 22151
rect 21315 22148 21327 22151
rect 21450 22148 21456 22160
rect 21315 22120 21456 22148
rect 21315 22117 21327 22120
rect 21269 22111 21327 22117
rect 21450 22108 21456 22120
rect 21508 22148 21514 22160
rect 21508 22120 21956 22148
rect 21508 22108 21514 22120
rect 17957 22083 18015 22089
rect 17957 22080 17969 22083
rect 17788 22052 17969 22080
rect 17674 22043 17732 22049
rect 17957 22049 17969 22052
rect 18003 22080 18015 22083
rect 18966 22080 18972 22092
rect 18003 22052 18972 22080
rect 18003 22049 18015 22052
rect 17957 22043 18015 22049
rect 14737 22015 14795 22021
rect 14016 21984 14228 22012
rect 13630 21944 13636 21956
rect 11388 21916 12112 21944
rect 12636 21916 13636 21944
rect 11388 21904 11394 21916
rect 12636 21888 12664 21916
rect 13630 21904 13636 21916
rect 13688 21904 13694 21956
rect 14200 21944 14228 21984
rect 14737 21981 14749 22015
rect 14783 22012 14795 22015
rect 15010 22012 15016 22024
rect 14783 21984 15016 22012
rect 14783 21981 14795 21984
rect 14737 21975 14795 21981
rect 15010 21972 15016 21984
rect 15068 21972 15074 22024
rect 15105 22015 15163 22021
rect 15105 21981 15117 22015
rect 15151 22012 15163 22015
rect 15470 22012 15476 22024
rect 15151 21984 15476 22012
rect 15151 21981 15163 21984
rect 15105 21975 15163 21981
rect 15470 21972 15476 21984
rect 15528 21972 15534 22024
rect 16482 21972 16488 22024
rect 16540 22012 16546 22024
rect 17512 22012 17540 22043
rect 18966 22040 18972 22052
rect 19024 22040 19030 22092
rect 19061 22083 19119 22089
rect 19061 22049 19073 22083
rect 19107 22080 19119 22083
rect 19150 22080 19156 22092
rect 19107 22052 19156 22080
rect 19107 22049 19119 22052
rect 19061 22043 19119 22049
rect 19150 22040 19156 22052
rect 19208 22040 19214 22092
rect 19702 22040 19708 22092
rect 19760 22040 19766 22092
rect 19794 22040 19800 22092
rect 19852 22080 19858 22092
rect 19981 22083 20039 22089
rect 19981 22080 19993 22083
rect 19852 22052 19993 22080
rect 19852 22040 19858 22052
rect 19981 22049 19993 22052
rect 20027 22049 20039 22083
rect 19981 22043 20039 22049
rect 20901 22083 20959 22089
rect 20901 22049 20913 22083
rect 20947 22080 20959 22083
rect 20990 22080 20996 22092
rect 20947 22052 20996 22080
rect 20947 22049 20959 22052
rect 20901 22043 20959 22049
rect 20990 22040 20996 22052
rect 21048 22040 21054 22092
rect 21361 22083 21419 22089
rect 21361 22049 21373 22083
rect 21407 22049 21419 22083
rect 21361 22043 21419 22049
rect 16540 21984 17540 22012
rect 16540 21972 16546 21984
rect 17586 21972 17592 22024
rect 17644 21972 17650 22024
rect 18049 22015 18107 22021
rect 18049 21981 18061 22015
rect 18095 22012 18107 22015
rect 18138 22012 18144 22024
rect 18095 21984 18144 22012
rect 18095 21981 18107 21984
rect 18049 21975 18107 21981
rect 18138 21972 18144 21984
rect 18196 22012 18202 22024
rect 19242 22012 19248 22024
rect 18196 21984 19248 22012
rect 18196 21972 18202 21984
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 21376 22012 21404 22043
rect 21542 22040 21548 22092
rect 21600 22040 21606 22092
rect 21634 22040 21640 22092
rect 21692 22040 21698 22092
rect 21928 22089 21956 22120
rect 22296 22089 22324 22188
rect 22554 22108 22560 22160
rect 22612 22108 22618 22160
rect 21913 22083 21971 22089
rect 21913 22080 21925 22083
rect 21891 22052 21925 22080
rect 21913 22049 21925 22052
rect 21959 22049 21971 22083
rect 21913 22043 21971 22049
rect 22281 22083 22339 22089
rect 22281 22049 22293 22083
rect 22327 22080 22339 22083
rect 22373 22083 22431 22089
rect 22373 22080 22385 22083
rect 22327 22052 22385 22080
rect 22327 22049 22339 22052
rect 22281 22043 22339 22049
rect 22373 22049 22385 22052
rect 22419 22049 22431 22083
rect 22373 22043 22431 22049
rect 21376 21984 21588 22012
rect 21560 21956 21588 21984
rect 15194 21944 15200 21956
rect 14200 21916 15200 21944
rect 15194 21904 15200 21916
rect 15252 21904 15258 21956
rect 21174 21944 21180 21956
rect 17788 21916 21180 21944
rect 9398 21876 9404 21888
rect 6420 21848 9404 21876
rect 6420 21836 6426 21848
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 11885 21879 11943 21885
rect 11885 21845 11897 21879
rect 11931 21876 11943 21879
rect 12618 21876 12624 21888
rect 11931 21848 12624 21876
rect 11931 21845 11943 21848
rect 11885 21839 11943 21845
rect 12618 21836 12624 21848
rect 12676 21836 12682 21888
rect 12897 21879 12955 21885
rect 12897 21845 12909 21879
rect 12943 21876 12955 21879
rect 12986 21876 12992 21888
rect 12943 21848 12992 21876
rect 12943 21845 12955 21848
rect 12897 21839 12955 21845
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 14826 21836 14832 21888
rect 14884 21836 14890 21888
rect 15470 21836 15476 21888
rect 15528 21876 15534 21888
rect 17788 21876 17816 21916
rect 15528 21848 17816 21876
rect 15528 21836 15534 21848
rect 17954 21836 17960 21888
rect 18012 21876 18018 21888
rect 19260 21885 19288 21916
rect 21174 21904 21180 21916
rect 21232 21904 21238 21956
rect 21542 21904 21548 21956
rect 21600 21904 21606 21956
rect 21652 21944 21680 22040
rect 21818 21972 21824 22024
rect 21876 22012 21882 22024
rect 22005 22015 22063 22021
rect 22005 22012 22017 22015
rect 21876 21984 22017 22012
rect 21876 21972 21882 21984
rect 22005 21981 22017 21984
rect 22051 21981 22063 22015
rect 22005 21975 22063 21981
rect 22186 21972 22192 22024
rect 22244 22012 22250 22024
rect 22741 22015 22799 22021
rect 22741 22012 22753 22015
rect 22244 21984 22753 22012
rect 22244 21972 22250 21984
rect 22741 21981 22753 21984
rect 22787 21981 22799 22015
rect 22741 21975 22799 21981
rect 21910 21944 21916 21956
rect 21652 21916 21916 21944
rect 21910 21904 21916 21916
rect 21968 21944 21974 21956
rect 21968 21916 22232 21944
rect 21968 21904 21974 21916
rect 18601 21879 18659 21885
rect 18601 21876 18613 21879
rect 18012 21848 18613 21876
rect 18012 21836 18018 21848
rect 18601 21845 18613 21848
rect 18647 21845 18659 21879
rect 18601 21839 18659 21845
rect 19245 21879 19303 21885
rect 19245 21845 19257 21879
rect 19291 21845 19303 21879
rect 19245 21839 19303 21845
rect 19794 21836 19800 21888
rect 19852 21876 19858 21888
rect 20533 21879 20591 21885
rect 20533 21876 20545 21879
rect 19852 21848 20545 21876
rect 19852 21836 19858 21848
rect 20533 21845 20545 21848
rect 20579 21876 20591 21879
rect 20622 21876 20628 21888
rect 20579 21848 20628 21876
rect 20579 21845 20591 21848
rect 20533 21839 20591 21845
rect 20622 21836 20628 21848
rect 20680 21836 20686 21888
rect 21726 21836 21732 21888
rect 21784 21836 21790 21888
rect 22094 21836 22100 21888
rect 22152 21836 22158 21888
rect 22204 21885 22232 21916
rect 22189 21879 22247 21885
rect 22189 21845 22201 21879
rect 22235 21845 22247 21879
rect 22189 21839 22247 21845
rect 552 21786 23368 21808
rect 552 21734 3662 21786
rect 3714 21734 3726 21786
rect 3778 21734 3790 21786
rect 3842 21734 3854 21786
rect 3906 21734 3918 21786
rect 3970 21734 23368 21786
rect 552 21712 23368 21734
rect 9030 21632 9036 21684
rect 9088 21672 9094 21684
rect 9398 21672 9404 21684
rect 9088 21644 9404 21672
rect 9088 21632 9094 21644
rect 9398 21632 9404 21644
rect 9456 21672 9462 21684
rect 9456 21644 10088 21672
rect 9456 21632 9462 21644
rect 4706 21564 4712 21616
rect 4764 21604 4770 21616
rect 5258 21604 5264 21616
rect 4764 21576 5264 21604
rect 4764 21564 4770 21576
rect 5258 21564 5264 21576
rect 5316 21564 5322 21616
rect 6273 21607 6331 21613
rect 6273 21573 6285 21607
rect 6319 21604 6331 21607
rect 7558 21604 7564 21616
rect 6319 21576 7564 21604
rect 6319 21573 6331 21576
rect 6273 21567 6331 21573
rect 7558 21564 7564 21576
rect 7616 21564 7622 21616
rect 8113 21607 8171 21613
rect 8113 21573 8125 21607
rect 8159 21604 8171 21607
rect 9585 21607 9643 21613
rect 8159 21576 9260 21604
rect 8159 21573 8171 21576
rect 8113 21567 8171 21573
rect 9232 21548 9260 21576
rect 9585 21573 9597 21607
rect 9631 21604 9643 21607
rect 9858 21604 9864 21616
rect 9631 21576 9864 21604
rect 9631 21573 9643 21576
rect 9585 21567 9643 21573
rect 9858 21564 9864 21576
rect 9916 21564 9922 21616
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21536 6055 21539
rect 6178 21536 6184 21548
rect 6043 21508 6184 21536
rect 6043 21505 6055 21508
rect 5997 21499 6055 21505
rect 6178 21496 6184 21508
rect 6236 21496 6242 21548
rect 6362 21496 6368 21548
rect 6420 21496 6426 21548
rect 7190 21496 7196 21548
rect 7248 21496 7254 21548
rect 7466 21496 7472 21548
rect 7524 21536 7530 21548
rect 7653 21539 7711 21545
rect 7653 21536 7665 21539
rect 7524 21508 7665 21536
rect 7524 21496 7530 21508
rect 7653 21505 7665 21508
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 8478 21496 8484 21548
rect 8536 21536 8542 21548
rect 8849 21539 8907 21545
rect 8849 21536 8861 21539
rect 8536 21508 8861 21536
rect 8536 21496 8542 21508
rect 8849 21505 8861 21508
rect 8895 21505 8907 21539
rect 8849 21499 8907 21505
rect 9033 21539 9091 21545
rect 9033 21505 9045 21539
rect 9079 21505 9091 21539
rect 9033 21499 9091 21505
rect 5905 21471 5963 21477
rect 5905 21437 5917 21471
rect 5951 21468 5963 21471
rect 6380 21468 6408 21496
rect 5951 21440 6408 21468
rect 5951 21437 5963 21440
rect 5905 21431 5963 21437
rect 4985 21403 5043 21409
rect 4985 21369 4997 21403
rect 5031 21400 5043 21403
rect 5074 21400 5080 21412
rect 5031 21372 5080 21400
rect 5031 21369 5043 21372
rect 4985 21363 5043 21369
rect 5074 21360 5080 21372
rect 5132 21400 5138 21412
rect 5258 21400 5264 21412
rect 5132 21372 5264 21400
rect 5132 21360 5138 21372
rect 5258 21360 5264 21372
rect 5316 21360 5322 21412
rect 6362 21360 6368 21412
rect 6420 21360 6426 21412
rect 7300 21400 7328 21454
rect 7742 21428 7748 21480
rect 7800 21428 7806 21480
rect 8570 21428 8576 21480
rect 8628 21468 8634 21480
rect 9048 21468 9076 21499
rect 9214 21496 9220 21548
rect 9272 21496 9278 21548
rect 9677 21539 9735 21545
rect 9677 21505 9689 21539
rect 9723 21536 9735 21539
rect 9723 21508 9996 21536
rect 9723 21505 9735 21508
rect 9677 21499 9735 21505
rect 9582 21468 9588 21480
rect 8628 21440 9588 21468
rect 8628 21428 8634 21440
rect 9582 21428 9588 21440
rect 9640 21428 9646 21480
rect 9766 21428 9772 21480
rect 9824 21428 9830 21480
rect 7650 21400 7656 21412
rect 7300 21372 7656 21400
rect 7650 21360 7656 21372
rect 7708 21400 7714 21412
rect 8110 21400 8116 21412
rect 7708 21372 8116 21400
rect 7708 21360 7714 21372
rect 8110 21360 8116 21372
rect 8168 21360 8174 21412
rect 8202 21360 8208 21412
rect 8260 21400 8266 21412
rect 8757 21403 8815 21409
rect 8757 21400 8769 21403
rect 8260 21372 8769 21400
rect 8260 21360 8266 21372
rect 8757 21369 8769 21372
rect 8803 21400 8815 21403
rect 9784 21400 9812 21428
rect 8803 21372 9812 21400
rect 9968 21400 9996 21508
rect 10060 21477 10088 21644
rect 12158 21632 12164 21684
rect 12216 21672 12222 21684
rect 13078 21672 13084 21684
rect 12216 21644 13084 21672
rect 12216 21632 12222 21644
rect 13078 21632 13084 21644
rect 13136 21632 13142 21684
rect 13446 21632 13452 21684
rect 13504 21672 13510 21684
rect 16761 21675 16819 21681
rect 13504 21644 13860 21672
rect 13504 21632 13510 21644
rect 10229 21607 10287 21613
rect 10229 21573 10241 21607
rect 10275 21604 10287 21607
rect 10275 21576 10824 21604
rect 10275 21573 10287 21576
rect 10229 21567 10287 21573
rect 10796 21536 10824 21576
rect 10870 21564 10876 21616
rect 10928 21564 10934 21616
rect 12618 21564 12624 21616
rect 12676 21604 12682 21616
rect 12676 21576 13124 21604
rect 12676 21564 12682 21576
rect 11974 21536 11980 21548
rect 10152 21508 10732 21536
rect 10796 21508 11980 21536
rect 10045 21471 10103 21477
rect 10045 21437 10057 21471
rect 10091 21437 10103 21471
rect 10045 21431 10103 21437
rect 10152 21400 10180 21508
rect 10226 21428 10232 21480
rect 10284 21468 10290 21480
rect 10704 21477 10732 21508
rect 11974 21496 11980 21508
rect 12032 21496 12038 21548
rect 12066 21496 12072 21548
rect 12124 21496 12130 21548
rect 12250 21496 12256 21548
rect 12308 21536 12314 21548
rect 12308 21508 12388 21536
rect 12308 21496 12314 21508
rect 10413 21471 10471 21477
rect 10413 21468 10425 21471
rect 10284 21440 10425 21468
rect 10284 21428 10290 21440
rect 10413 21437 10425 21440
rect 10459 21437 10471 21471
rect 10413 21431 10471 21437
rect 10689 21471 10747 21477
rect 10689 21437 10701 21471
rect 10735 21437 10747 21471
rect 10689 21431 10747 21437
rect 9968 21372 10180 21400
rect 10428 21400 10456 21431
rect 10778 21428 10784 21480
rect 10836 21468 10842 21480
rect 11057 21471 11115 21477
rect 11057 21468 11069 21471
rect 10836 21440 11069 21468
rect 10836 21428 10842 21440
rect 11057 21437 11069 21440
rect 11103 21437 11115 21471
rect 12360 21468 12388 21508
rect 12436 21471 12494 21477
rect 12436 21468 12448 21471
rect 11057 21431 11115 21437
rect 10428 21372 10916 21400
rect 8803 21369 8815 21372
rect 8757 21363 8815 21369
rect 5166 21292 5172 21344
rect 5224 21332 5230 21344
rect 5445 21335 5503 21341
rect 5445 21332 5457 21335
rect 5224 21304 5457 21332
rect 5224 21292 5230 21304
rect 5445 21301 5457 21304
rect 5491 21301 5503 21335
rect 5445 21295 5503 21301
rect 8389 21335 8447 21341
rect 8389 21301 8401 21335
rect 8435 21332 8447 21335
rect 8478 21332 8484 21344
rect 8435 21304 8484 21332
rect 8435 21301 8447 21304
rect 8389 21295 8447 21301
rect 8478 21292 8484 21304
rect 8536 21292 8542 21344
rect 9766 21292 9772 21344
rect 9824 21332 9830 21344
rect 9861 21335 9919 21341
rect 9861 21332 9873 21335
rect 9824 21304 9873 21332
rect 9824 21292 9830 21304
rect 9861 21301 9873 21304
rect 9907 21301 9919 21335
rect 9861 21295 9919 21301
rect 10505 21335 10563 21341
rect 10505 21301 10517 21335
rect 10551 21332 10563 21335
rect 10778 21332 10784 21344
rect 10551 21304 10784 21332
rect 10551 21301 10563 21304
rect 10505 21295 10563 21301
rect 10778 21292 10784 21304
rect 10836 21292 10842 21344
rect 10888 21332 10916 21372
rect 11164 21332 11192 21454
rect 12360 21440 12448 21468
rect 12436 21437 12448 21440
rect 12482 21437 12494 21471
rect 12436 21431 12494 21437
rect 12529 21471 12587 21477
rect 12529 21437 12541 21471
rect 12575 21468 12587 21471
rect 12802 21468 12808 21480
rect 12575 21440 12808 21468
rect 12575 21437 12587 21440
rect 12529 21431 12587 21437
rect 12802 21428 12808 21440
rect 12860 21428 12866 21480
rect 13096 21477 13124 21576
rect 13262 21564 13268 21616
rect 13320 21604 13326 21616
rect 13357 21607 13415 21613
rect 13357 21604 13369 21607
rect 13320 21576 13369 21604
rect 13320 21564 13326 21576
rect 13357 21573 13369 21576
rect 13403 21604 13415 21607
rect 13722 21604 13728 21616
rect 13403 21576 13728 21604
rect 13403 21573 13415 21576
rect 13357 21567 13415 21573
rect 13722 21564 13728 21576
rect 13780 21564 13786 21616
rect 13832 21604 13860 21644
rect 16761 21641 16773 21675
rect 16807 21672 16819 21675
rect 17218 21672 17224 21684
rect 16807 21644 17224 21672
rect 16807 21641 16819 21644
rect 16761 21635 16819 21641
rect 17218 21632 17224 21644
rect 17276 21672 17282 21684
rect 17770 21672 17776 21684
rect 17276 21644 17776 21672
rect 17276 21632 17282 21644
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 19794 21672 19800 21684
rect 18156 21644 19800 21672
rect 15565 21607 15623 21613
rect 15565 21604 15577 21607
rect 13832 21576 15577 21604
rect 15565 21573 15577 21576
rect 15611 21573 15623 21607
rect 17313 21607 17371 21613
rect 17313 21604 17325 21607
rect 15565 21567 15623 21573
rect 16592 21576 17325 21604
rect 13538 21536 13544 21548
rect 13188 21508 13544 21536
rect 13188 21477 13216 21508
rect 13538 21496 13544 21508
rect 13596 21496 13602 21548
rect 14642 21496 14648 21548
rect 14700 21496 14706 21548
rect 16592 21545 16620 21576
rect 17313 21573 17325 21576
rect 17359 21573 17371 21607
rect 17313 21567 17371 21573
rect 17402 21564 17408 21616
rect 17460 21604 17466 21616
rect 18156 21604 18184 21644
rect 19794 21632 19800 21644
rect 19852 21632 19858 21684
rect 21450 21632 21456 21684
rect 21508 21632 21514 21684
rect 22186 21672 22192 21684
rect 21836 21644 22192 21672
rect 17460 21576 18184 21604
rect 18233 21607 18291 21613
rect 17460 21564 17466 21576
rect 18233 21573 18245 21607
rect 18279 21604 18291 21607
rect 18874 21604 18880 21616
rect 18279 21576 18880 21604
rect 18279 21573 18291 21576
rect 18233 21567 18291 21573
rect 18874 21564 18880 21576
rect 18932 21604 18938 21616
rect 21836 21613 21864 21644
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 19613 21607 19671 21613
rect 18932 21576 19452 21604
rect 18932 21564 18938 21576
rect 16025 21539 16083 21545
rect 16025 21505 16037 21539
rect 16071 21536 16083 21539
rect 16577 21539 16635 21545
rect 16577 21536 16589 21539
rect 16071 21508 16589 21536
rect 16071 21505 16083 21508
rect 16025 21499 16083 21505
rect 16577 21505 16589 21508
rect 16623 21505 16635 21539
rect 16577 21499 16635 21505
rect 17034 21496 17040 21548
rect 17092 21536 17098 21548
rect 18414 21536 18420 21548
rect 17092 21508 18420 21536
rect 17092 21496 17098 21508
rect 13081 21471 13139 21477
rect 13081 21437 13093 21471
rect 13127 21437 13139 21471
rect 13081 21431 13139 21437
rect 13173 21471 13231 21477
rect 13173 21437 13185 21471
rect 13219 21437 13231 21471
rect 13173 21431 13231 21437
rect 13354 21428 13360 21480
rect 13412 21428 13418 21480
rect 13909 21471 13967 21477
rect 13909 21437 13921 21471
rect 13955 21437 13967 21471
rect 13909 21431 13967 21437
rect 12342 21360 12348 21412
rect 12400 21400 12406 21412
rect 12710 21400 12716 21412
rect 12400 21372 12716 21400
rect 12400 21360 12406 21372
rect 12710 21360 12716 21372
rect 12768 21360 12774 21412
rect 13924 21400 13952 21431
rect 13998 21428 14004 21480
rect 14056 21468 14062 21480
rect 14458 21468 14464 21480
rect 14056 21440 14464 21468
rect 14056 21428 14062 21440
rect 14458 21428 14464 21440
rect 14516 21428 14522 21480
rect 14734 21428 14740 21480
rect 14792 21428 14798 21480
rect 15930 21428 15936 21480
rect 15988 21428 15994 21480
rect 16390 21428 16396 21480
rect 16448 21468 16454 21480
rect 16485 21471 16543 21477
rect 16485 21468 16497 21471
rect 16448 21440 16497 21468
rect 16448 21428 16454 21440
rect 16485 21437 16497 21440
rect 16531 21468 16543 21471
rect 16531 21440 17080 21468
rect 16531 21437 16543 21440
rect 16485 21431 16543 21437
rect 14752 21400 14780 21428
rect 13924 21372 14780 21400
rect 16114 21360 16120 21412
rect 16172 21400 16178 21412
rect 16945 21403 17003 21409
rect 16945 21400 16957 21403
rect 16172 21372 16957 21400
rect 16172 21360 16178 21372
rect 16945 21369 16957 21372
rect 16991 21369 17003 21403
rect 17052 21400 17080 21440
rect 17126 21428 17132 21480
rect 17184 21428 17190 21480
rect 17310 21428 17316 21480
rect 17368 21468 17374 21480
rect 17681 21471 17739 21477
rect 17681 21468 17693 21471
rect 17368 21440 17693 21468
rect 17368 21428 17374 21440
rect 17681 21437 17693 21440
rect 17727 21437 17739 21471
rect 17681 21431 17739 21437
rect 17865 21471 17923 21477
rect 17865 21437 17877 21471
rect 17911 21468 17923 21471
rect 17954 21468 17960 21480
rect 17911 21440 17960 21468
rect 17911 21437 17923 21440
rect 17865 21431 17923 21437
rect 17954 21428 17960 21440
rect 18012 21428 18018 21480
rect 18064 21477 18092 21508
rect 18414 21496 18420 21508
rect 18472 21496 18478 21548
rect 18969 21539 19027 21545
rect 18969 21536 18981 21539
rect 18708 21508 18981 21536
rect 18049 21471 18107 21477
rect 18049 21437 18061 21471
rect 18095 21437 18107 21471
rect 18049 21431 18107 21437
rect 18230 21428 18236 21480
rect 18288 21428 18294 21480
rect 18509 21471 18567 21477
rect 18509 21437 18521 21471
rect 18555 21462 18567 21471
rect 18708 21468 18736 21508
rect 18969 21505 18981 21508
rect 19015 21536 19027 21539
rect 19058 21536 19064 21548
rect 19015 21508 19064 21536
rect 19015 21505 19027 21508
rect 18969 21499 19027 21505
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 19242 21496 19248 21548
rect 19300 21496 19306 21548
rect 18632 21462 18736 21468
rect 18555 21440 18736 21462
rect 18555 21437 18660 21440
rect 18509 21434 18660 21437
rect 18509 21431 18567 21434
rect 18874 21428 18880 21480
rect 18932 21428 18938 21480
rect 19337 21471 19395 21477
rect 19337 21437 19349 21471
rect 19383 21437 19395 21471
rect 19337 21431 19395 21437
rect 17402 21400 17408 21412
rect 17052 21372 17408 21400
rect 16945 21363 17003 21369
rect 17402 21360 17408 21372
rect 17460 21360 17466 21412
rect 18417 21403 18475 21409
rect 18417 21369 18429 21403
rect 18463 21400 18475 21403
rect 19352 21400 19380 21431
rect 18463 21372 19380 21400
rect 19424 21400 19452 21576
rect 19613 21573 19625 21607
rect 19659 21573 19671 21607
rect 19613 21567 19671 21573
rect 21821 21607 21879 21613
rect 21821 21573 21833 21607
rect 21867 21573 21879 21607
rect 22097 21607 22155 21613
rect 22097 21604 22109 21607
rect 21821 21567 21879 21573
rect 21928 21576 22109 21604
rect 19628 21468 19656 21567
rect 21928 21536 21956 21576
rect 22097 21573 22109 21576
rect 22143 21573 22155 21607
rect 22097 21567 22155 21573
rect 20732 21508 21956 21536
rect 22005 21539 22063 21545
rect 20732 21480 20760 21508
rect 22005 21505 22017 21539
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 20530 21468 20536 21480
rect 20588 21477 20594 21480
rect 20588 21471 20621 21477
rect 19628 21440 20536 21468
rect 20530 21428 20536 21440
rect 20609 21437 20621 21471
rect 20588 21431 20621 21437
rect 20588 21428 20594 21431
rect 20714 21428 20720 21480
rect 20772 21428 20778 21480
rect 20990 21428 20996 21480
rect 21048 21428 21054 21480
rect 21082 21428 21088 21480
rect 21140 21428 21146 21480
rect 21269 21471 21327 21477
rect 21269 21437 21281 21471
rect 21315 21468 21327 21471
rect 21358 21468 21364 21480
rect 21315 21440 21364 21468
rect 21315 21437 21327 21440
rect 21269 21431 21327 21437
rect 21358 21428 21364 21440
rect 21416 21428 21422 21480
rect 22020 21468 22048 21499
rect 22097 21471 22155 21477
rect 22097 21468 22109 21471
rect 22020 21440 22109 21468
rect 22097 21437 22109 21440
rect 22143 21437 22155 21471
rect 22097 21431 22155 21437
rect 22281 21471 22339 21477
rect 22281 21437 22293 21471
rect 22327 21437 22339 21471
rect 22281 21431 22339 21437
rect 19613 21403 19671 21409
rect 19613 21400 19625 21403
rect 19424 21372 19625 21400
rect 18463 21369 18475 21372
rect 18417 21363 18475 21369
rect 19613 21369 19625 21372
rect 19659 21369 19671 21403
rect 19613 21363 19671 21369
rect 21174 21360 21180 21412
rect 21232 21400 21238 21412
rect 21545 21403 21603 21409
rect 21545 21400 21557 21403
rect 21232 21372 21557 21400
rect 21232 21360 21238 21372
rect 21545 21369 21557 21372
rect 21591 21369 21603 21403
rect 21545 21363 21603 21369
rect 10888 21304 11192 21332
rect 12158 21292 12164 21344
rect 12216 21292 12222 21344
rect 13541 21335 13599 21341
rect 13541 21301 13553 21335
rect 13587 21332 13599 21335
rect 14090 21332 14096 21344
rect 13587 21304 14096 21332
rect 13587 21301 13599 21304
rect 13541 21295 13599 21301
rect 14090 21292 14096 21304
rect 14148 21292 14154 21344
rect 14182 21292 14188 21344
rect 14240 21292 14246 21344
rect 15286 21292 15292 21344
rect 15344 21332 15350 21344
rect 15381 21335 15439 21341
rect 15381 21332 15393 21335
rect 15344 21304 15393 21332
rect 15344 21292 15350 21304
rect 15381 21301 15393 21304
rect 15427 21301 15439 21335
rect 15381 21295 15439 21301
rect 17494 21292 17500 21344
rect 17552 21292 17558 21344
rect 18874 21292 18880 21344
rect 18932 21332 18938 21344
rect 19429 21335 19487 21341
rect 19429 21332 19441 21335
rect 18932 21304 19441 21332
rect 18932 21292 18938 21304
rect 19429 21301 19441 21304
rect 19475 21301 19487 21335
rect 19429 21295 19487 21301
rect 20349 21335 20407 21341
rect 20349 21301 20361 21335
rect 20395 21332 20407 21335
rect 20438 21332 20444 21344
rect 20395 21304 20444 21332
rect 20395 21301 20407 21304
rect 20349 21295 20407 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 21560 21332 21588 21363
rect 21910 21360 21916 21412
rect 21968 21400 21974 21412
rect 22296 21400 22324 21431
rect 21968 21372 22324 21400
rect 21968 21360 21974 21372
rect 22002 21332 22008 21344
rect 21560 21304 22008 21332
rect 22002 21292 22008 21304
rect 22060 21292 22066 21344
rect 552 21242 23368 21264
rect 552 21190 4322 21242
rect 4374 21190 4386 21242
rect 4438 21190 4450 21242
rect 4502 21190 4514 21242
rect 4566 21190 4578 21242
rect 4630 21190 23368 21242
rect 552 21168 23368 21190
rect 5626 21088 5632 21140
rect 5684 21128 5690 21140
rect 6362 21128 6368 21140
rect 5684 21100 6368 21128
rect 5684 21088 5690 21100
rect 6362 21088 6368 21100
rect 6420 21128 6426 21140
rect 6420 21100 6500 21128
rect 6420 21088 6426 21100
rect 5166 21020 5172 21072
rect 5224 21060 5230 21072
rect 6472 21069 6500 21100
rect 8110 21088 8116 21140
rect 8168 21128 8174 21140
rect 9766 21128 9772 21140
rect 8168 21100 9772 21128
rect 8168 21088 8174 21100
rect 7932 21072 7984 21078
rect 6457 21063 6515 21069
rect 5224 21032 6224 21060
rect 5224 21020 5230 21032
rect 4525 20995 4583 21001
rect 4525 20961 4537 20995
rect 4571 20992 4583 20995
rect 4985 20995 5043 21001
rect 4985 20992 4997 20995
rect 4571 20964 4997 20992
rect 4571 20961 4583 20964
rect 4525 20955 4583 20961
rect 4985 20961 4997 20964
rect 5031 20992 5043 20995
rect 5258 20992 5264 21004
rect 5031 20964 5264 20992
rect 5031 20961 5043 20964
rect 4985 20955 5043 20961
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 5626 20952 5632 21004
rect 5684 20992 5690 21004
rect 6196 21001 6224 21032
rect 6457 21029 6469 21063
rect 6503 21029 6515 21063
rect 6457 21023 6515 21029
rect 7932 21014 7984 21020
rect 5905 20995 5963 21001
rect 5905 20992 5917 20995
rect 5684 20964 5917 20992
rect 5684 20952 5690 20964
rect 5905 20961 5917 20964
rect 5951 20961 5963 20995
rect 5905 20955 5963 20961
rect 6181 20995 6239 21001
rect 6181 20961 6193 20995
rect 6227 20961 6239 20995
rect 6181 20955 6239 20961
rect 6641 20995 6699 21001
rect 6641 20961 6653 20995
rect 6687 20992 6699 20995
rect 6914 20992 6920 21004
rect 6687 20964 6920 20992
rect 6687 20961 6699 20964
rect 6641 20955 6699 20961
rect 6914 20952 6920 20964
rect 6972 20992 6978 21004
rect 7098 20992 7104 21004
rect 6972 20964 7104 20992
rect 6972 20952 6978 20964
rect 7098 20952 7104 20964
rect 7156 20952 7162 21004
rect 8202 20952 8208 21004
rect 8260 20952 8266 21004
rect 8849 20995 8907 21001
rect 8849 20961 8861 20995
rect 8895 20992 8907 20995
rect 8956 20992 8984 21100
rect 9766 21088 9772 21100
rect 9824 21128 9830 21140
rect 10689 21131 10747 21137
rect 9824 21100 10548 21128
rect 9824 21088 9830 21100
rect 9398 21020 9404 21072
rect 9456 21060 9462 21072
rect 10229 21063 10287 21069
rect 9456 21032 10180 21060
rect 9456 21020 9462 21032
rect 8895 20964 8984 20992
rect 8895 20961 8907 20964
rect 8849 20955 8907 20961
rect 9490 20952 9496 21004
rect 9548 20952 9554 21004
rect 9674 20952 9680 21004
rect 9732 20952 9738 21004
rect 9769 20995 9827 21001
rect 9769 20961 9781 20995
rect 9815 20992 9827 20995
rect 9950 20992 9956 21004
rect 9815 20964 9956 20992
rect 9815 20961 9827 20964
rect 9769 20955 9827 20961
rect 9950 20952 9956 20964
rect 10008 20952 10014 21004
rect 10152 21001 10180 21032
rect 10229 21029 10241 21063
rect 10275 21060 10287 21063
rect 10520 21060 10548 21100
rect 10689 21097 10701 21131
rect 10735 21128 10747 21131
rect 10778 21128 10784 21140
rect 10735 21100 10784 21128
rect 10735 21097 10747 21100
rect 10689 21091 10747 21097
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 11241 21131 11299 21137
rect 11241 21097 11253 21131
rect 11287 21128 11299 21131
rect 11698 21128 11704 21140
rect 11287 21100 11704 21128
rect 11287 21097 11299 21100
rect 11241 21091 11299 21097
rect 11698 21088 11704 21100
rect 11756 21088 11762 21140
rect 12342 21128 12348 21140
rect 11808 21100 12348 21128
rect 11808 21060 11836 21100
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 14090 21088 14096 21140
rect 14148 21088 14154 21140
rect 16482 21088 16488 21140
rect 16540 21088 16546 21140
rect 17310 21088 17316 21140
rect 17368 21088 17374 21140
rect 14737 21063 14795 21069
rect 10275 21032 10456 21060
rect 10520 21032 11836 21060
rect 12406 21032 14688 21060
rect 10275 21029 10287 21032
rect 10229 21023 10287 21029
rect 10137 20995 10195 21001
rect 10137 20961 10149 20995
rect 10183 20961 10195 20995
rect 10137 20955 10195 20961
rect 10318 20952 10324 21004
rect 10376 20952 10382 21004
rect 10428 20992 10456 21032
rect 10597 20995 10655 21001
rect 10597 20992 10609 20995
rect 10428 20964 10609 20992
rect 10597 20961 10609 20964
rect 10643 20961 10655 20995
rect 10597 20955 10655 20961
rect 10778 20952 10784 21004
rect 10836 20952 10842 21004
rect 11054 20952 11060 21004
rect 11112 20952 11118 21004
rect 11422 20952 11428 21004
rect 11480 20992 11486 21004
rect 12406 20992 12434 21032
rect 11480 20964 12434 20992
rect 11480 20952 11486 20964
rect 13170 20952 13176 21004
rect 13228 20992 13234 21004
rect 13725 20995 13783 21001
rect 13725 20992 13737 20995
rect 13228 20964 13737 20992
rect 13228 20952 13234 20964
rect 13725 20961 13737 20964
rect 13771 20961 13783 20995
rect 13725 20955 13783 20961
rect 13906 20952 13912 21004
rect 13964 20952 13970 21004
rect 4614 20884 4620 20936
rect 4672 20884 4678 20936
rect 4709 20927 4767 20933
rect 4709 20893 4721 20927
rect 4755 20893 4767 20927
rect 4709 20887 4767 20893
rect 4724 20856 4752 20887
rect 5074 20884 5080 20936
rect 5132 20924 5138 20936
rect 6089 20927 6147 20933
rect 6089 20924 6101 20927
rect 5132 20896 6101 20924
rect 5132 20884 5138 20896
rect 6089 20893 6101 20896
rect 6135 20893 6147 20927
rect 11606 20924 11612 20936
rect 6089 20887 6147 20893
rect 9646 20896 11612 20924
rect 5350 20856 5356 20868
rect 4724 20828 5356 20856
rect 5350 20816 5356 20828
rect 5408 20816 5414 20868
rect 5997 20859 6055 20865
rect 5997 20825 6009 20859
rect 6043 20825 6055 20859
rect 5997 20819 6055 20825
rect 6365 20859 6423 20865
rect 6365 20825 6377 20859
rect 6411 20856 6423 20859
rect 9646 20856 9674 20896
rect 11606 20884 11612 20896
rect 11664 20884 11670 20936
rect 14660 20924 14688 21032
rect 14737 21029 14749 21063
rect 14783 21060 14795 21063
rect 14918 21060 14924 21072
rect 14783 21032 14924 21060
rect 14783 21029 14795 21032
rect 14737 21023 14795 21029
rect 14918 21020 14924 21032
rect 14976 21020 14982 21072
rect 15930 21020 15936 21072
rect 15988 21060 15994 21072
rect 20990 21060 20996 21072
rect 15988 21032 20996 21060
rect 15988 21020 15994 21032
rect 20990 21020 20996 21032
rect 21048 21020 21054 21072
rect 15010 20952 15016 21004
rect 15068 20952 15074 21004
rect 15470 20952 15476 21004
rect 15528 20952 15534 21004
rect 16298 20952 16304 21004
rect 16356 20952 16362 21004
rect 16485 20995 16543 21001
rect 16485 20961 16497 20995
rect 16531 20961 16543 20995
rect 16485 20955 16543 20961
rect 15746 20924 15752 20936
rect 14660 20896 15752 20924
rect 15746 20884 15752 20896
rect 15804 20924 15810 20936
rect 16500 20924 16528 20955
rect 17218 20952 17224 21004
rect 17276 20952 17282 21004
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20992 17463 20995
rect 17586 20992 17592 21004
rect 17451 20964 17592 20992
rect 17451 20961 17463 20964
rect 17405 20955 17463 20961
rect 17586 20952 17592 20964
rect 17644 20952 17650 21004
rect 20257 20995 20315 21001
rect 20257 20961 20269 20995
rect 20303 20961 20315 20995
rect 20257 20955 20315 20961
rect 15804 20896 16528 20924
rect 20272 20924 20300 20955
rect 20438 20952 20444 21004
rect 20496 20952 20502 21004
rect 20530 20952 20536 21004
rect 20588 20952 20594 21004
rect 20714 21001 20720 21004
rect 20687 20995 20720 21001
rect 20687 20961 20699 20995
rect 20687 20955 20720 20961
rect 20714 20952 20720 20955
rect 20772 20952 20778 21004
rect 20901 20995 20959 21001
rect 20901 20961 20913 20995
rect 20947 20992 20959 20995
rect 21082 20992 21088 21004
rect 20947 20964 21088 20992
rect 20947 20961 20959 20964
rect 20901 20955 20959 20961
rect 20916 20924 20944 20955
rect 21082 20952 21088 20964
rect 21140 20992 21146 21004
rect 21637 20995 21695 21001
rect 21637 20992 21649 20995
rect 21140 20964 21649 20992
rect 21140 20952 21146 20964
rect 21637 20961 21649 20964
rect 21683 20961 21695 20995
rect 21637 20955 21695 20961
rect 21726 20952 21732 21004
rect 21784 20992 21790 21004
rect 22373 20995 22431 21001
rect 22373 20992 22385 20995
rect 21784 20964 22385 20992
rect 21784 20952 21790 20964
rect 22373 20961 22385 20964
rect 22419 20961 22431 20995
rect 22373 20955 22431 20961
rect 20272 20896 20944 20924
rect 21453 20927 21511 20933
rect 15804 20884 15810 20896
rect 21453 20893 21465 20927
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 6411 20828 9674 20856
rect 6411 20825 6423 20828
rect 6365 20819 6423 20825
rect 4893 20791 4951 20797
rect 4893 20757 4905 20791
rect 4939 20788 4951 20791
rect 5074 20788 5080 20800
rect 4939 20760 5080 20788
rect 4939 20757 4951 20760
rect 4893 20751 4951 20757
rect 5074 20748 5080 20760
rect 5132 20748 5138 20800
rect 5442 20748 5448 20800
rect 5500 20788 5506 20800
rect 6012 20788 6040 20819
rect 10318 20816 10324 20868
rect 10376 20856 10382 20868
rect 15930 20856 15936 20868
rect 10376 20828 15936 20856
rect 10376 20816 10382 20828
rect 15930 20816 15936 20828
rect 15988 20816 15994 20868
rect 21468 20856 21496 20887
rect 21542 20884 21548 20936
rect 21600 20884 21606 20936
rect 22094 20856 22100 20868
rect 21468 20828 22100 20856
rect 22094 20816 22100 20828
rect 22152 20816 22158 20868
rect 5500 20760 6040 20788
rect 5500 20748 5506 20760
rect 6638 20748 6644 20800
rect 6696 20788 6702 20800
rect 6825 20791 6883 20797
rect 6825 20788 6837 20791
rect 6696 20760 6837 20788
rect 6696 20748 6702 20760
rect 6825 20757 6837 20760
rect 6871 20757 6883 20791
rect 6825 20751 6883 20757
rect 9122 20748 9128 20800
rect 9180 20788 9186 20800
rect 9309 20791 9367 20797
rect 9309 20788 9321 20791
rect 9180 20760 9321 20788
rect 9180 20748 9186 20760
rect 9309 20757 9321 20760
rect 9355 20757 9367 20791
rect 9309 20751 9367 20757
rect 9490 20748 9496 20800
rect 9548 20788 9554 20800
rect 11146 20788 11152 20800
rect 9548 20760 11152 20788
rect 9548 20748 9554 20760
rect 11146 20748 11152 20760
rect 11204 20748 11210 20800
rect 11330 20748 11336 20800
rect 11388 20788 11394 20800
rect 11425 20791 11483 20797
rect 11425 20788 11437 20791
rect 11388 20760 11437 20788
rect 11388 20748 11394 20760
rect 11425 20757 11437 20760
rect 11471 20757 11483 20791
rect 11425 20751 11483 20757
rect 13722 20748 13728 20800
rect 13780 20748 13786 20800
rect 20254 20748 20260 20800
rect 20312 20788 20318 20800
rect 20349 20791 20407 20797
rect 20349 20788 20361 20791
rect 20312 20760 20361 20788
rect 20312 20748 20318 20760
rect 20349 20757 20361 20760
rect 20395 20757 20407 20791
rect 20349 20751 20407 20757
rect 21266 20748 21272 20800
rect 21324 20748 21330 20800
rect 21910 20748 21916 20800
rect 21968 20748 21974 20800
rect 552 20698 23368 20720
rect 552 20646 3662 20698
rect 3714 20646 3726 20698
rect 3778 20646 3790 20698
rect 3842 20646 3854 20698
rect 3906 20646 3918 20698
rect 3970 20646 23368 20698
rect 552 20624 23368 20646
rect 5074 20544 5080 20596
rect 5132 20544 5138 20596
rect 5442 20544 5448 20596
rect 5500 20584 5506 20596
rect 5997 20587 6055 20593
rect 5997 20584 6009 20587
rect 5500 20556 6009 20584
rect 5500 20544 5506 20556
rect 5997 20553 6009 20556
rect 6043 20553 6055 20587
rect 5997 20547 6055 20553
rect 6086 20544 6092 20596
rect 6144 20584 6150 20596
rect 8662 20584 8668 20596
rect 6144 20556 8668 20584
rect 6144 20544 6150 20556
rect 8662 20544 8668 20556
rect 8720 20584 8726 20596
rect 10134 20584 10140 20596
rect 8720 20556 10140 20584
rect 8720 20544 8726 20556
rect 10134 20544 10140 20556
rect 10192 20544 10198 20596
rect 10321 20587 10379 20593
rect 10321 20553 10333 20587
rect 10367 20584 10379 20587
rect 10778 20584 10784 20596
rect 10367 20556 10784 20584
rect 10367 20553 10379 20556
rect 10321 20547 10379 20553
rect 10778 20544 10784 20556
rect 10836 20584 10842 20596
rect 13170 20584 13176 20596
rect 10836 20556 13176 20584
rect 10836 20544 10842 20556
rect 13170 20544 13176 20556
rect 13228 20584 13234 20596
rect 13228 20556 13584 20584
rect 13228 20544 13234 20556
rect 5092 20516 5120 20544
rect 7009 20519 7067 20525
rect 5092 20488 6132 20516
rect 5166 20408 5172 20460
rect 5224 20408 5230 20460
rect 5626 20408 5632 20460
rect 5684 20408 5690 20460
rect 5902 20408 5908 20460
rect 5960 20408 5966 20460
rect 6104 20457 6132 20488
rect 7009 20485 7021 20519
rect 7055 20516 7067 20519
rect 7055 20488 13492 20516
rect 7055 20485 7067 20488
rect 7009 20479 7067 20485
rect 6089 20451 6147 20457
rect 6089 20417 6101 20451
rect 6135 20417 6147 20451
rect 7024 20448 7052 20479
rect 6089 20411 6147 20417
rect 6840 20420 7052 20448
rect 5261 20383 5319 20389
rect 5261 20349 5273 20383
rect 5307 20380 5319 20383
rect 5442 20380 5448 20392
rect 5307 20352 5448 20380
rect 5307 20349 5319 20352
rect 5261 20343 5319 20349
rect 5442 20340 5448 20352
rect 5500 20340 5506 20392
rect 5537 20383 5595 20389
rect 5537 20349 5549 20383
rect 5583 20349 5595 20383
rect 5537 20343 5595 20349
rect 4893 20247 4951 20253
rect 4893 20213 4905 20247
rect 4939 20244 4951 20247
rect 5552 20244 5580 20343
rect 5644 20312 5672 20408
rect 5994 20340 6000 20392
rect 6052 20340 6058 20392
rect 6638 20340 6644 20392
rect 6696 20340 6702 20392
rect 6840 20389 6868 20420
rect 10870 20408 10876 20460
rect 10928 20448 10934 20460
rect 12342 20448 12348 20460
rect 10928 20420 12348 20448
rect 10928 20408 10934 20420
rect 12342 20408 12348 20420
rect 12400 20448 12406 20460
rect 12400 20420 12848 20448
rect 12400 20408 12406 20420
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 6917 20383 6975 20389
rect 6917 20349 6929 20383
rect 6963 20349 6975 20383
rect 6917 20343 6975 20349
rect 6932 20312 6960 20343
rect 7098 20340 7104 20392
rect 7156 20340 7162 20392
rect 7926 20340 7932 20392
rect 7984 20380 7990 20392
rect 8389 20383 8447 20389
rect 8389 20380 8401 20383
rect 7984 20352 8401 20380
rect 7984 20340 7990 20352
rect 8389 20349 8401 20352
rect 8435 20349 8447 20383
rect 8389 20343 8447 20349
rect 8481 20383 8539 20389
rect 8481 20349 8493 20383
rect 8527 20380 8539 20383
rect 8570 20380 8576 20392
rect 8527 20352 8576 20380
rect 8527 20349 8539 20352
rect 8481 20343 8539 20349
rect 8570 20340 8576 20352
rect 8628 20340 8634 20392
rect 8662 20340 8668 20392
rect 8720 20340 8726 20392
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 10042 20380 10048 20392
rect 9732 20352 10048 20380
rect 9732 20340 9738 20352
rect 10042 20340 10048 20352
rect 10100 20380 10106 20392
rect 10321 20383 10379 20389
rect 10321 20380 10333 20383
rect 10100 20352 10333 20380
rect 10100 20340 10106 20352
rect 10321 20349 10333 20352
rect 10367 20349 10379 20383
rect 10321 20343 10379 20349
rect 10505 20383 10563 20389
rect 10505 20349 10517 20383
rect 10551 20380 10563 20383
rect 10962 20380 10968 20392
rect 10551 20352 10968 20380
rect 10551 20349 10563 20352
rect 10505 20343 10563 20349
rect 10962 20340 10968 20352
rect 11020 20340 11026 20392
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 12820 20389 12848 20420
rect 12621 20383 12679 20389
rect 12621 20380 12633 20383
rect 12492 20352 12633 20380
rect 12492 20340 12498 20352
rect 12621 20349 12633 20352
rect 12667 20349 12679 20383
rect 12621 20343 12679 20349
rect 12805 20383 12863 20389
rect 12805 20349 12817 20383
rect 12851 20349 12863 20383
rect 13464 20380 13492 20488
rect 13556 20457 13584 20556
rect 14642 20544 14648 20596
rect 14700 20544 14706 20596
rect 21269 20587 21327 20593
rect 21269 20584 21281 20587
rect 20732 20556 21281 20584
rect 15562 20516 15568 20528
rect 13648 20488 15568 20516
rect 13541 20451 13599 20457
rect 13541 20417 13553 20451
rect 13587 20417 13599 20451
rect 13541 20411 13599 20417
rect 13648 20380 13676 20488
rect 15562 20476 15568 20488
rect 15620 20516 15626 20528
rect 16298 20516 16304 20528
rect 15620 20488 16304 20516
rect 15620 20476 15626 20488
rect 16298 20476 16304 20488
rect 16356 20476 16362 20528
rect 14090 20408 14096 20460
rect 14148 20448 14154 20460
rect 14277 20451 14335 20457
rect 14277 20448 14289 20451
rect 14148 20420 14289 20448
rect 14148 20408 14154 20420
rect 14277 20417 14289 20420
rect 14323 20417 14335 20451
rect 14277 20411 14335 20417
rect 14366 20408 14372 20460
rect 14424 20448 14430 20460
rect 16390 20448 16396 20460
rect 14424 20420 16396 20448
rect 14424 20408 14430 20420
rect 16390 20408 16396 20420
rect 16448 20408 16454 20460
rect 17221 20451 17279 20457
rect 17221 20417 17233 20451
rect 17267 20417 17279 20451
rect 17221 20411 17279 20417
rect 17512 20420 17724 20448
rect 13464 20352 13676 20380
rect 12805 20343 12863 20349
rect 13722 20340 13728 20392
rect 13780 20340 13786 20392
rect 14458 20340 14464 20392
rect 14516 20340 14522 20392
rect 5644 20284 6960 20312
rect 7374 20272 7380 20324
rect 7432 20312 7438 20324
rect 17236 20312 17264 20411
rect 17512 20392 17540 20420
rect 17313 20383 17371 20389
rect 17313 20349 17325 20383
rect 17359 20380 17371 20383
rect 17494 20380 17500 20392
rect 17359 20352 17500 20380
rect 17359 20349 17371 20352
rect 17313 20343 17371 20349
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 17696 20389 17724 20420
rect 20732 20392 20760 20556
rect 21269 20553 21281 20556
rect 21315 20584 21327 20587
rect 21542 20584 21548 20596
rect 21315 20556 21548 20584
rect 21315 20553 21327 20556
rect 21269 20547 21327 20553
rect 21542 20544 21548 20556
rect 21600 20544 21606 20596
rect 20993 20519 21051 20525
rect 20993 20485 21005 20519
rect 21039 20516 21051 20519
rect 22646 20516 22652 20528
rect 21039 20488 22652 20516
rect 21039 20485 21051 20488
rect 20993 20479 21051 20485
rect 22646 20476 22652 20488
rect 22704 20476 22710 20528
rect 17589 20383 17647 20389
rect 17589 20349 17601 20383
rect 17635 20349 17647 20383
rect 17589 20343 17647 20349
rect 17682 20383 17740 20389
rect 17682 20349 17694 20383
rect 17728 20349 17740 20383
rect 17682 20343 17740 20349
rect 17604 20312 17632 20343
rect 18322 20340 18328 20392
rect 18380 20380 18386 20392
rect 18693 20383 18751 20389
rect 18693 20380 18705 20383
rect 18380 20352 18705 20380
rect 18380 20340 18386 20352
rect 18693 20349 18705 20352
rect 18739 20349 18751 20383
rect 18693 20343 18751 20349
rect 18874 20340 18880 20392
rect 18932 20340 18938 20392
rect 20530 20340 20536 20392
rect 20588 20380 20594 20392
rect 20625 20383 20683 20389
rect 20625 20380 20637 20383
rect 20588 20352 20637 20380
rect 20588 20340 20594 20352
rect 20625 20349 20637 20352
rect 20671 20349 20683 20383
rect 20625 20343 20683 20349
rect 7432 20284 17632 20312
rect 7432 20272 7438 20284
rect 5718 20244 5724 20256
rect 4939 20216 5724 20244
rect 4939 20213 4951 20216
rect 4893 20207 4951 20213
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 6362 20204 6368 20256
rect 6420 20204 6426 20256
rect 6825 20247 6883 20253
rect 6825 20213 6837 20247
rect 6871 20244 6883 20247
rect 6914 20244 6920 20256
rect 6871 20216 6920 20244
rect 6871 20213 6883 20216
rect 6825 20207 6883 20213
rect 6914 20204 6920 20216
rect 6972 20204 6978 20256
rect 8849 20247 8907 20253
rect 8849 20213 8861 20247
rect 8895 20244 8907 20247
rect 8938 20244 8944 20256
rect 8895 20216 8944 20244
rect 8895 20213 8907 20216
rect 8849 20207 8907 20213
rect 8938 20204 8944 20216
rect 8996 20204 9002 20256
rect 12989 20247 13047 20253
rect 12989 20213 13001 20247
rect 13035 20244 13047 20247
rect 13630 20244 13636 20256
rect 13035 20216 13636 20244
rect 13035 20213 13047 20216
rect 12989 20207 13047 20213
rect 13630 20204 13636 20216
rect 13688 20204 13694 20256
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 13909 20247 13967 20253
rect 13909 20244 13921 20247
rect 13872 20216 13921 20244
rect 13872 20204 13878 20216
rect 13909 20213 13921 20216
rect 13955 20213 13967 20247
rect 13909 20207 13967 20213
rect 16945 20247 17003 20253
rect 16945 20213 16957 20247
rect 16991 20244 17003 20247
rect 17126 20244 17132 20256
rect 16991 20216 17132 20244
rect 16991 20213 17003 20216
rect 16945 20207 17003 20213
rect 17126 20204 17132 20216
rect 17184 20204 17190 20256
rect 17957 20247 18015 20253
rect 17957 20213 17969 20247
rect 18003 20244 18015 20247
rect 18138 20244 18144 20256
rect 18003 20216 18144 20244
rect 18003 20213 18015 20216
rect 17957 20207 18015 20213
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 18506 20204 18512 20256
rect 18564 20244 18570 20256
rect 18785 20247 18843 20253
rect 18785 20244 18797 20247
rect 18564 20216 18797 20244
rect 18564 20204 18570 20216
rect 18785 20213 18797 20216
rect 18831 20213 18843 20247
rect 18785 20207 18843 20213
rect 20438 20204 20444 20256
rect 20496 20204 20502 20256
rect 20640 20244 20668 20343
rect 20714 20340 20720 20392
rect 20772 20340 20778 20392
rect 20993 20383 21051 20389
rect 20993 20349 21005 20383
rect 21039 20380 21051 20383
rect 21910 20380 21916 20392
rect 21039 20352 21916 20380
rect 21039 20349 21051 20352
rect 20993 20343 21051 20349
rect 20809 20315 20867 20321
rect 20809 20281 20821 20315
rect 20855 20312 20867 20315
rect 21082 20312 21088 20324
rect 20855 20284 21088 20312
rect 20855 20281 20867 20284
rect 20809 20275 20867 20281
rect 21082 20272 21088 20284
rect 21140 20272 21146 20324
rect 21284 20321 21312 20352
rect 21910 20340 21916 20352
rect 21968 20340 21974 20392
rect 22186 20340 22192 20392
rect 22244 20340 22250 20392
rect 21284 20315 21343 20321
rect 21284 20284 21297 20315
rect 21285 20281 21297 20284
rect 21331 20281 21343 20315
rect 21285 20275 21343 20281
rect 21376 20284 21588 20312
rect 21376 20244 21404 20284
rect 20640 20216 21404 20244
rect 21450 20204 21456 20256
rect 21508 20204 21514 20256
rect 21560 20244 21588 20284
rect 21634 20272 21640 20324
rect 21692 20312 21698 20324
rect 21729 20315 21787 20321
rect 21729 20312 21741 20315
rect 21692 20284 21741 20312
rect 21692 20272 21698 20284
rect 21729 20281 21741 20284
rect 21775 20281 21787 20315
rect 21729 20275 21787 20281
rect 21821 20247 21879 20253
rect 21821 20244 21833 20247
rect 21560 20216 21833 20244
rect 21821 20213 21833 20216
rect 21867 20213 21879 20247
rect 21821 20207 21879 20213
rect 22370 20204 22376 20256
rect 22428 20204 22434 20256
rect 552 20154 23368 20176
rect 552 20102 4322 20154
rect 4374 20102 4386 20154
rect 4438 20102 4450 20154
rect 4502 20102 4514 20154
rect 4566 20102 4578 20154
rect 4630 20102 23368 20154
rect 552 20080 23368 20102
rect 7374 20000 7380 20052
rect 7432 20000 7438 20052
rect 7926 20040 7932 20052
rect 7484 20012 7932 20040
rect 5994 19932 6000 19984
rect 6052 19972 6058 19984
rect 7484 19972 7512 20012
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 11701 20043 11759 20049
rect 11701 20009 11713 20043
rect 11747 20040 11759 20043
rect 13541 20043 13599 20049
rect 11747 20012 12434 20040
rect 11747 20009 11759 20012
rect 11701 20003 11759 20009
rect 8570 19972 8576 19984
rect 6052 19944 7512 19972
rect 7852 19944 8576 19972
rect 6052 19932 6058 19944
rect 5534 19864 5540 19916
rect 5592 19904 5598 19916
rect 5905 19907 5963 19913
rect 5905 19904 5917 19907
rect 5592 19876 5917 19904
rect 5592 19864 5598 19876
rect 5905 19873 5917 19876
rect 5951 19873 5963 19907
rect 5905 19867 5963 19873
rect 6086 19864 6092 19916
rect 6144 19904 6150 19916
rect 6181 19907 6239 19913
rect 6181 19904 6193 19907
rect 6144 19876 6193 19904
rect 6144 19864 6150 19876
rect 6181 19873 6193 19876
rect 6227 19873 6239 19907
rect 6181 19867 6239 19873
rect 6641 19907 6699 19913
rect 6641 19873 6653 19907
rect 6687 19904 6699 19907
rect 6914 19904 6920 19916
rect 6687 19876 6920 19904
rect 6687 19873 6699 19876
rect 6641 19867 6699 19873
rect 6914 19864 6920 19876
rect 6972 19864 6978 19916
rect 7558 19864 7564 19916
rect 7616 19864 7622 19916
rect 7852 19913 7880 19944
rect 8570 19932 8576 19944
rect 8628 19972 8634 19984
rect 8849 19975 8907 19981
rect 8849 19972 8861 19975
rect 8628 19944 8861 19972
rect 8628 19932 8634 19944
rect 8849 19941 8861 19944
rect 8895 19941 8907 19975
rect 8849 19935 8907 19941
rect 12406 19916 12434 20012
rect 13541 20009 13553 20043
rect 13587 20040 13599 20043
rect 13587 20012 14228 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 13630 19932 13636 19984
rect 13688 19932 13694 19984
rect 7837 19907 7895 19913
rect 7837 19873 7849 19907
rect 7883 19873 7895 19907
rect 7837 19867 7895 19873
rect 8389 19907 8447 19913
rect 8389 19873 8401 19907
rect 8435 19904 8447 19907
rect 9766 19904 9772 19916
rect 8435 19876 9772 19904
rect 8435 19873 8447 19876
rect 8389 19867 8447 19873
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 10318 19864 10324 19916
rect 10376 19864 10382 19916
rect 10689 19907 10747 19913
rect 10689 19873 10701 19907
rect 10735 19904 10747 19907
rect 11054 19904 11060 19916
rect 10735 19876 11060 19904
rect 10735 19873 10747 19876
rect 10689 19867 10747 19873
rect 11054 19864 11060 19876
rect 11112 19904 11118 19916
rect 11333 19907 11391 19913
rect 11333 19904 11345 19907
rect 11112 19876 11345 19904
rect 11112 19864 11118 19876
rect 11333 19873 11345 19876
rect 11379 19873 11391 19907
rect 12406 19876 12440 19916
rect 11333 19867 11391 19873
rect 12434 19864 12440 19876
rect 12492 19864 12498 19916
rect 13170 19864 13176 19916
rect 13228 19864 13234 19916
rect 13814 19864 13820 19916
rect 13872 19864 13878 19916
rect 13906 19864 13912 19916
rect 13964 19864 13970 19916
rect 14090 19864 14096 19916
rect 14148 19904 14154 19916
rect 14200 19913 14228 20012
rect 18138 20000 18144 20052
rect 18196 20000 18202 20052
rect 18414 20000 18420 20052
rect 18472 20040 18478 20052
rect 18782 20040 18788 20052
rect 18472 20012 18788 20040
rect 18472 20000 18478 20012
rect 18782 20000 18788 20012
rect 18840 20040 18846 20052
rect 19242 20049 19248 20052
rect 19229 20043 19248 20049
rect 19229 20040 19241 20043
rect 18840 20012 19241 20040
rect 18840 20000 18846 20012
rect 19229 20009 19241 20012
rect 19229 20003 19248 20009
rect 19242 20000 19248 20003
rect 19300 20000 19306 20052
rect 20165 20043 20223 20049
rect 20165 20009 20177 20043
rect 20211 20040 20223 20043
rect 20346 20040 20352 20052
rect 20211 20012 20352 20040
rect 20211 20009 20223 20012
rect 20165 20003 20223 20009
rect 20346 20000 20352 20012
rect 20404 20040 20410 20052
rect 20714 20040 20720 20052
rect 20404 20012 20720 20040
rect 20404 20000 20410 20012
rect 20714 20000 20720 20012
rect 20772 20000 20778 20052
rect 21266 20000 21272 20052
rect 21324 20000 21330 20052
rect 21450 20000 21456 20052
rect 21508 20040 21514 20052
rect 21508 20012 22508 20040
rect 21508 20000 21514 20012
rect 17037 19975 17095 19981
rect 17037 19941 17049 19975
rect 17083 19972 17095 19975
rect 18156 19972 18184 20000
rect 19429 19975 19487 19981
rect 17083 19944 18092 19972
rect 18156 19944 18644 19972
rect 17083 19941 17095 19944
rect 17037 19935 17095 19941
rect 14185 19907 14243 19913
rect 14185 19904 14197 19907
rect 14148 19876 14197 19904
rect 14148 19864 14154 19876
rect 14185 19873 14197 19876
rect 14231 19873 14243 19907
rect 14185 19867 14243 19873
rect 16390 19864 16396 19916
rect 16448 19904 16454 19916
rect 16945 19907 17003 19913
rect 16945 19904 16957 19907
rect 16448 19876 16957 19904
rect 16448 19864 16454 19876
rect 16945 19873 16957 19876
rect 16991 19873 17003 19907
rect 16945 19867 17003 19873
rect 6549 19839 6607 19845
rect 6549 19805 6561 19839
rect 6595 19805 6607 19839
rect 6549 19799 6607 19805
rect 6181 19771 6239 19777
rect 6181 19737 6193 19771
rect 6227 19768 6239 19771
rect 6564 19768 6592 19799
rect 8294 19796 8300 19848
rect 8352 19796 8358 19848
rect 11238 19796 11244 19848
rect 11296 19796 11302 19848
rect 12342 19796 12348 19848
rect 12400 19796 12406 19848
rect 12805 19839 12863 19845
rect 12805 19805 12817 19839
rect 12851 19836 12863 19839
rect 13265 19839 13323 19845
rect 13265 19836 13277 19839
rect 12851 19808 13277 19836
rect 12851 19805 12863 19808
rect 12805 19799 12863 19805
rect 13265 19805 13277 19808
rect 13311 19836 13323 19839
rect 13722 19836 13728 19848
rect 13311 19808 13728 19836
rect 13311 19805 13323 19808
rect 13265 19799 13323 19805
rect 13722 19796 13728 19808
rect 13780 19796 13786 19848
rect 14274 19796 14280 19848
rect 14332 19836 14338 19848
rect 14826 19836 14832 19848
rect 14332 19808 14832 19836
rect 14332 19796 14338 19808
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 6822 19768 6828 19780
rect 6227 19740 6828 19768
rect 6227 19737 6239 19740
rect 6181 19731 6239 19737
rect 6822 19728 6828 19740
rect 6880 19728 6886 19780
rect 7009 19771 7067 19777
rect 7009 19737 7021 19771
rect 7055 19768 7067 19771
rect 7742 19768 7748 19780
rect 7055 19740 7748 19768
rect 7055 19737 7067 19740
rect 7009 19731 7067 19737
rect 7742 19728 7748 19740
rect 7800 19728 7806 19780
rect 8757 19771 8815 19777
rect 8757 19737 8769 19771
rect 8803 19768 8815 19771
rect 9490 19768 9496 19780
rect 8803 19740 9496 19768
rect 8803 19737 8815 19740
rect 8757 19731 8815 19737
rect 9490 19728 9496 19740
rect 9548 19728 9554 19780
rect 13909 19771 13967 19777
rect 13909 19737 13921 19771
rect 13955 19768 13967 19771
rect 14734 19768 14740 19780
rect 13955 19740 14740 19768
rect 13955 19737 13967 19740
rect 13909 19731 13967 19737
rect 14734 19728 14740 19740
rect 14792 19728 14798 19780
rect 16960 19768 16988 19867
rect 17126 19864 17132 19916
rect 17184 19904 17190 19916
rect 18064 19913 18092 19944
rect 17405 19907 17463 19913
rect 17184 19876 17356 19904
rect 17184 19864 17190 19876
rect 17328 19845 17356 19876
rect 17405 19873 17417 19907
rect 17451 19873 17463 19907
rect 17405 19867 17463 19873
rect 18049 19907 18107 19913
rect 18049 19873 18061 19907
rect 18095 19873 18107 19907
rect 18049 19867 18107 19873
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18414 19904 18420 19916
rect 18371 19876 18420 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 17313 19839 17371 19845
rect 17313 19805 17325 19839
rect 17359 19805 17371 19839
rect 17313 19799 17371 19805
rect 17420 19768 17448 19867
rect 18064 19836 18092 19867
rect 18414 19864 18420 19876
rect 18472 19864 18478 19916
rect 18506 19864 18512 19916
rect 18564 19864 18570 19916
rect 18616 19913 18644 19944
rect 19429 19941 19441 19975
rect 19475 19941 19487 19975
rect 21284 19972 21312 20000
rect 19429 19935 19487 19941
rect 19812 19944 20392 19972
rect 18601 19907 18659 19913
rect 18601 19873 18613 19907
rect 18647 19904 18659 19907
rect 19444 19904 19472 19935
rect 19812 19916 19840 19944
rect 18647 19876 19472 19904
rect 19705 19907 19763 19913
rect 18647 19873 18659 19876
rect 18601 19867 18659 19873
rect 19705 19873 19717 19907
rect 19751 19873 19763 19907
rect 19705 19867 19763 19873
rect 18693 19839 18751 19845
rect 18693 19836 18705 19839
rect 18064 19808 18705 19836
rect 16960 19740 17448 19768
rect 17773 19771 17831 19777
rect 17773 19737 17785 19771
rect 17819 19768 17831 19771
rect 17954 19768 17960 19780
rect 17819 19740 17960 19768
rect 17819 19737 17831 19740
rect 17773 19731 17831 19737
rect 17954 19728 17960 19740
rect 18012 19728 18018 19780
rect 10962 19660 10968 19712
rect 11020 19700 11026 19712
rect 14366 19700 14372 19712
rect 11020 19672 14372 19700
rect 11020 19660 11026 19672
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 14553 19703 14611 19709
rect 14553 19669 14565 19703
rect 14599 19700 14611 19703
rect 15102 19700 15108 19712
rect 14599 19672 15108 19700
rect 14599 19669 14611 19672
rect 14553 19663 14611 19669
rect 15102 19660 15108 19672
rect 15160 19660 15166 19712
rect 18248 19700 18276 19808
rect 18693 19805 18705 19808
rect 18739 19805 18751 19839
rect 18693 19799 18751 19805
rect 18782 19796 18788 19848
rect 18840 19796 18846 19848
rect 18969 19839 19027 19845
rect 18969 19805 18981 19839
rect 19015 19836 19027 19839
rect 19720 19836 19748 19867
rect 19794 19864 19800 19916
rect 19852 19864 19858 19916
rect 19981 19907 20039 19913
rect 19981 19873 19993 19907
rect 20027 19904 20039 19907
rect 20254 19904 20260 19916
rect 20027 19876 20260 19904
rect 20027 19873 20039 19876
rect 19981 19867 20039 19873
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 20364 19913 20392 19944
rect 20732 19944 21312 19972
rect 21913 19975 21971 19981
rect 20349 19907 20407 19913
rect 20349 19873 20361 19907
rect 20395 19873 20407 19907
rect 20349 19867 20407 19873
rect 20533 19907 20591 19913
rect 20533 19873 20545 19907
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 20548 19836 20576 19867
rect 20622 19864 20628 19916
rect 20680 19864 20686 19916
rect 20732 19913 20760 19944
rect 21913 19941 21925 19975
rect 21959 19972 21971 19975
rect 22189 19975 22247 19981
rect 22189 19972 22201 19975
rect 21959 19944 22201 19972
rect 21959 19941 21971 19944
rect 21913 19935 21971 19941
rect 22189 19941 22201 19944
rect 22235 19941 22247 19975
rect 22189 19935 22247 19941
rect 20717 19907 20775 19913
rect 20717 19873 20729 19907
rect 20763 19873 20775 19907
rect 20717 19867 20775 19873
rect 20901 19907 20959 19913
rect 20901 19873 20913 19907
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 19015 19808 20576 19836
rect 19015 19805 19027 19808
rect 18969 19799 19027 19805
rect 18322 19728 18328 19780
rect 18380 19728 18386 19780
rect 18984 19740 19288 19768
rect 18984 19700 19012 19740
rect 18248 19672 19012 19700
rect 19058 19660 19064 19712
rect 19116 19660 19122 19712
rect 19260 19709 19288 19740
rect 20622 19728 20628 19780
rect 20680 19768 20686 19780
rect 20916 19768 20944 19867
rect 21082 19864 21088 19916
rect 21140 19904 21146 19916
rect 22005 19907 22063 19913
rect 22005 19904 22017 19907
rect 21140 19876 22017 19904
rect 21140 19864 21146 19876
rect 22005 19873 22017 19876
rect 22051 19873 22063 19907
rect 22005 19867 22063 19873
rect 22278 19864 22284 19916
rect 22336 19864 22342 19916
rect 22370 19864 22376 19916
rect 22428 19864 22434 19916
rect 22480 19904 22508 20012
rect 22649 19907 22707 19913
rect 22649 19904 22661 19907
rect 22480 19876 22661 19904
rect 22649 19873 22661 19876
rect 22695 19873 22707 19907
rect 22649 19867 22707 19873
rect 20990 19796 20996 19848
rect 21048 19836 21054 19848
rect 21637 19839 21695 19845
rect 21637 19836 21649 19839
rect 21048 19808 21649 19836
rect 21048 19796 21054 19808
rect 21637 19805 21649 19808
rect 21683 19805 21695 19839
rect 21637 19799 21695 19805
rect 21726 19796 21732 19848
rect 21784 19796 21790 19848
rect 22388 19836 22416 19864
rect 22741 19839 22799 19845
rect 22741 19836 22753 19839
rect 22388 19808 22753 19836
rect 22741 19805 22753 19808
rect 22787 19805 22799 19839
rect 22741 19799 22799 19805
rect 20680 19740 20944 19768
rect 20680 19728 20686 19740
rect 19245 19703 19303 19709
rect 19245 19669 19257 19703
rect 19291 19669 19303 19703
rect 19245 19663 19303 19669
rect 20254 19660 20260 19712
rect 20312 19660 20318 19712
rect 22462 19660 22468 19712
rect 22520 19700 22526 19712
rect 22557 19703 22615 19709
rect 22557 19700 22569 19703
rect 22520 19672 22569 19700
rect 22520 19660 22526 19672
rect 22557 19669 22569 19672
rect 22603 19669 22615 19703
rect 22557 19663 22615 19669
rect 22646 19660 22652 19712
rect 22704 19660 22710 19712
rect 22738 19660 22744 19712
rect 22796 19700 22802 19712
rect 23017 19703 23075 19709
rect 23017 19700 23029 19703
rect 22796 19672 23029 19700
rect 22796 19660 22802 19672
rect 23017 19669 23029 19672
rect 23063 19669 23075 19703
rect 23017 19663 23075 19669
rect 552 19610 23368 19632
rect 552 19558 3662 19610
rect 3714 19558 3726 19610
rect 3778 19558 3790 19610
rect 3842 19558 3854 19610
rect 3906 19558 3918 19610
rect 3970 19558 23368 19610
rect 552 19536 23368 19558
rect 5626 19456 5632 19508
rect 5684 19456 5690 19508
rect 7193 19499 7251 19505
rect 7193 19465 7205 19499
rect 7239 19496 7251 19499
rect 7558 19496 7564 19508
rect 7239 19468 7564 19496
rect 7239 19465 7251 19468
rect 7193 19459 7251 19465
rect 7558 19456 7564 19468
rect 7616 19456 7622 19508
rect 8113 19499 8171 19505
rect 8113 19465 8125 19499
rect 8159 19496 8171 19499
rect 18509 19499 18567 19505
rect 8159 19468 15424 19496
rect 8159 19465 8171 19468
rect 8113 19459 8171 19465
rect 9585 19431 9643 19437
rect 9585 19397 9597 19431
rect 9631 19397 9643 19431
rect 9585 19391 9643 19397
rect 7742 19320 7748 19372
rect 7800 19320 7806 19372
rect 6822 19252 6828 19304
rect 6880 19252 6886 19304
rect 6914 19252 6920 19304
rect 6972 19292 6978 19304
rect 7009 19295 7067 19301
rect 7009 19292 7021 19295
rect 6972 19264 7021 19292
rect 6972 19252 6978 19264
rect 7009 19261 7021 19264
rect 7055 19261 7067 19295
rect 7009 19255 7067 19261
rect 7837 19295 7895 19301
rect 7837 19261 7849 19295
rect 7883 19261 7895 19295
rect 7837 19255 7895 19261
rect 4706 19184 4712 19236
rect 4764 19224 4770 19236
rect 5442 19224 5448 19236
rect 4764 19196 5448 19224
rect 4764 19184 4770 19196
rect 5442 19184 5448 19196
rect 5500 19184 5506 19236
rect 7558 19184 7564 19236
rect 7616 19224 7622 19236
rect 7852 19224 7880 19255
rect 8662 19252 8668 19304
rect 8720 19252 8726 19304
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19292 8907 19295
rect 9398 19292 9404 19304
rect 8895 19264 9404 19292
rect 8895 19261 8907 19264
rect 8849 19255 8907 19261
rect 9398 19252 9404 19264
rect 9456 19252 9462 19304
rect 9600 19224 9628 19391
rect 13630 19388 13636 19440
rect 13688 19388 13694 19440
rect 13541 19363 13599 19369
rect 13541 19329 13553 19363
rect 13587 19360 13599 19363
rect 13648 19360 13676 19388
rect 13587 19332 13676 19360
rect 14016 19332 14688 19360
rect 13587 19329 13599 19332
rect 13541 19323 13599 19329
rect 9769 19295 9827 19301
rect 9769 19261 9781 19295
rect 9815 19261 9827 19295
rect 9769 19255 9827 19261
rect 10413 19295 10471 19301
rect 10413 19261 10425 19295
rect 10459 19292 10471 19295
rect 10962 19292 10968 19304
rect 10459 19264 10968 19292
rect 10459 19261 10471 19264
rect 10413 19255 10471 19261
rect 9784 19224 9812 19255
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11974 19252 11980 19304
rect 12032 19252 12038 19304
rect 12805 19295 12863 19301
rect 12805 19261 12817 19295
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19292 13691 19295
rect 13722 19292 13728 19304
rect 13679 19264 13728 19292
rect 13679 19261 13691 19264
rect 13633 19255 13691 19261
rect 11054 19224 11060 19236
rect 7616 19196 9720 19224
rect 9784 19196 11060 19224
rect 7616 19184 7622 19196
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 5645 19159 5703 19165
rect 5645 19156 5657 19159
rect 5316 19128 5657 19156
rect 5316 19116 5322 19128
rect 5645 19125 5657 19128
rect 5691 19125 5703 19159
rect 5645 19119 5703 19125
rect 5813 19159 5871 19165
rect 5813 19125 5825 19159
rect 5859 19156 5871 19159
rect 7282 19156 7288 19168
rect 5859 19128 7288 19156
rect 5859 19125 5871 19128
rect 5813 19119 5871 19125
rect 7282 19116 7288 19128
rect 7340 19116 7346 19168
rect 8849 19159 8907 19165
rect 8849 19125 8861 19159
rect 8895 19156 8907 19159
rect 9582 19156 9588 19168
rect 8895 19128 9588 19156
rect 8895 19125 8907 19128
rect 8849 19119 8907 19125
rect 9582 19116 9588 19128
rect 9640 19116 9646 19168
rect 9692 19156 9720 19196
rect 11054 19184 11060 19196
rect 11112 19224 11118 19236
rect 11112 19196 11362 19224
rect 11112 19184 11118 19196
rect 12342 19184 12348 19236
rect 12400 19224 12406 19236
rect 12820 19224 12848 19255
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 13814 19252 13820 19304
rect 13872 19252 13878 19304
rect 14016 19292 14044 19332
rect 13924 19264 14044 19292
rect 13924 19224 13952 19264
rect 14090 19252 14096 19304
rect 14148 19252 14154 19304
rect 14274 19301 14280 19304
rect 14247 19295 14280 19301
rect 14247 19261 14259 19295
rect 14247 19255 14280 19261
rect 14274 19252 14280 19255
rect 14332 19252 14338 19304
rect 14550 19252 14556 19304
rect 14608 19252 14614 19304
rect 12400 19196 13952 19224
rect 14001 19227 14059 19233
rect 12400 19184 12406 19196
rect 14001 19193 14013 19227
rect 14047 19224 14059 19227
rect 14568 19224 14596 19252
rect 14047 19196 14596 19224
rect 14660 19224 14688 19332
rect 14734 19252 14740 19304
rect 14792 19252 14798 19304
rect 15396 19301 15424 19468
rect 18509 19465 18521 19499
rect 18555 19496 18567 19499
rect 18690 19496 18696 19508
rect 18555 19468 18696 19496
rect 18555 19465 18567 19468
rect 18509 19459 18567 19465
rect 18690 19456 18696 19468
rect 18748 19496 18754 19508
rect 18874 19496 18880 19508
rect 18748 19468 18880 19496
rect 18748 19456 18754 19468
rect 18874 19456 18880 19468
rect 18932 19456 18938 19508
rect 20717 19499 20775 19505
rect 20717 19465 20729 19499
rect 20763 19496 20775 19499
rect 22554 19496 22560 19508
rect 20763 19468 22560 19496
rect 20763 19465 20775 19468
rect 20717 19459 20775 19465
rect 22554 19456 22560 19468
rect 22612 19456 22618 19508
rect 16577 19431 16635 19437
rect 16577 19397 16589 19431
rect 16623 19397 16635 19431
rect 16577 19391 16635 19397
rect 15470 19320 15476 19372
rect 15528 19320 15534 19372
rect 15749 19363 15807 19369
rect 15749 19329 15761 19363
rect 15795 19360 15807 19363
rect 15795 19332 16344 19360
rect 15795 19329 15807 19332
rect 15749 19323 15807 19329
rect 16316 19304 16344 19332
rect 15381 19295 15439 19301
rect 15381 19261 15393 19295
rect 15427 19292 15439 19295
rect 15841 19295 15899 19301
rect 15841 19292 15853 19295
rect 15427 19264 15853 19292
rect 15427 19261 15439 19264
rect 15381 19255 15439 19261
rect 15841 19261 15853 19264
rect 15887 19261 15899 19295
rect 15841 19255 15899 19261
rect 16025 19295 16083 19301
rect 16025 19261 16037 19295
rect 16071 19261 16083 19295
rect 16025 19255 16083 19261
rect 14660 19196 15424 19224
rect 14047 19193 14059 19196
rect 14001 19187 14059 19193
rect 15396 19168 15424 19196
rect 15470 19184 15476 19236
rect 15528 19224 15534 19236
rect 16040 19224 16068 19255
rect 16298 19252 16304 19304
rect 16356 19252 16362 19304
rect 16390 19252 16396 19304
rect 16448 19252 16454 19304
rect 16592 19292 16620 19391
rect 18322 19388 18328 19440
rect 18380 19428 18386 19440
rect 18380 19400 18736 19428
rect 18380 19388 18386 19400
rect 17972 19332 18368 19360
rect 17972 19304 18000 19332
rect 16592 19264 17908 19292
rect 15528 19196 16068 19224
rect 16209 19227 16267 19233
rect 15528 19184 15534 19196
rect 16209 19193 16221 19227
rect 16255 19224 16267 19227
rect 16577 19227 16635 19233
rect 16577 19224 16589 19227
rect 16255 19196 16589 19224
rect 16255 19193 16267 19196
rect 16209 19187 16267 19193
rect 16577 19193 16589 19196
rect 16623 19193 16635 19227
rect 17880 19224 17908 19264
rect 17954 19252 17960 19304
rect 18012 19252 18018 19304
rect 18340 19301 18368 19332
rect 18708 19301 18736 19400
rect 20254 19388 20260 19440
rect 20312 19388 20318 19440
rect 20438 19388 20444 19440
rect 20496 19388 20502 19440
rect 20165 19363 20223 19369
rect 20165 19329 20177 19363
rect 20211 19360 20223 19363
rect 20272 19360 20300 19388
rect 20211 19332 20300 19360
rect 20349 19363 20407 19369
rect 20211 19329 20223 19332
rect 20165 19323 20223 19329
rect 20349 19329 20361 19363
rect 20395 19360 20407 19363
rect 20456 19360 20484 19388
rect 20395 19332 20484 19360
rect 20395 19329 20407 19332
rect 20349 19323 20407 19329
rect 18049 19295 18107 19301
rect 18049 19261 18061 19295
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18325 19295 18383 19301
rect 18325 19261 18337 19295
rect 18371 19261 18383 19295
rect 18325 19255 18383 19261
rect 18509 19295 18567 19301
rect 18509 19261 18521 19295
rect 18555 19261 18567 19295
rect 18509 19255 18567 19261
rect 18693 19295 18751 19301
rect 18693 19261 18705 19295
rect 18739 19261 18751 19295
rect 18693 19255 18751 19261
rect 18877 19295 18935 19301
rect 18877 19261 18889 19295
rect 18923 19292 18935 19295
rect 19058 19292 19064 19304
rect 18923 19264 19064 19292
rect 18923 19261 18935 19264
rect 18877 19255 18935 19261
rect 18064 19224 18092 19255
rect 18524 19224 18552 19255
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 20254 19252 20260 19304
rect 20312 19252 20318 19304
rect 17880 19196 18552 19224
rect 16577 19187 16635 19193
rect 19334 19184 19340 19236
rect 19392 19224 19398 19236
rect 20364 19224 20392 19323
rect 20438 19252 20444 19304
rect 20496 19252 20502 19304
rect 20622 19292 20628 19304
rect 20548 19264 20628 19292
rect 19392 19196 20392 19224
rect 19392 19184 19398 19196
rect 10134 19156 10140 19168
rect 9692 19128 10140 19156
rect 10134 19116 10140 19128
rect 10192 19116 10198 19168
rect 14458 19116 14464 19168
rect 14516 19116 14522 19168
rect 14645 19159 14703 19165
rect 14645 19125 14657 19159
rect 14691 19156 14703 19159
rect 14734 19156 14740 19168
rect 14691 19128 14740 19156
rect 14691 19125 14703 19128
rect 14645 19119 14703 19125
rect 14734 19116 14740 19128
rect 14792 19116 14798 19168
rect 15378 19116 15384 19168
rect 15436 19116 15442 19168
rect 18230 19116 18236 19168
rect 18288 19116 18294 19168
rect 18506 19116 18512 19168
rect 18564 19156 18570 19168
rect 18785 19159 18843 19165
rect 18785 19156 18797 19159
rect 18564 19128 18797 19156
rect 18564 19116 18570 19128
rect 18785 19125 18797 19128
rect 18831 19125 18843 19159
rect 18785 19119 18843 19125
rect 19978 19116 19984 19168
rect 20036 19116 20042 19168
rect 20162 19116 20168 19168
rect 20220 19156 20226 19168
rect 20548 19156 20576 19264
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 21082 19252 21088 19304
rect 21140 19292 21146 19304
rect 21140 19264 21185 19292
rect 21140 19252 21146 19264
rect 22462 19252 22468 19304
rect 22520 19301 22526 19304
rect 22520 19292 22532 19301
rect 22741 19295 22799 19301
rect 22520 19264 22565 19292
rect 22520 19255 22532 19264
rect 22741 19261 22753 19295
rect 22787 19292 22799 19295
rect 22830 19292 22836 19304
rect 22787 19264 22836 19292
rect 22787 19261 22799 19264
rect 22741 19255 22799 19261
rect 22520 19252 22526 19255
rect 22830 19252 22836 19264
rect 22888 19252 22894 19304
rect 21726 19224 21732 19236
rect 21100 19196 21732 19224
rect 21100 19165 21128 19196
rect 21726 19184 21732 19196
rect 21784 19184 21790 19236
rect 20220 19128 20576 19156
rect 21085 19159 21143 19165
rect 20220 19116 20226 19128
rect 21085 19125 21097 19159
rect 21131 19125 21143 19159
rect 21085 19119 21143 19125
rect 21266 19116 21272 19168
rect 21324 19116 21330 19168
rect 21361 19159 21419 19165
rect 21361 19125 21373 19159
rect 21407 19156 21419 19159
rect 22278 19156 22284 19168
rect 21407 19128 22284 19156
rect 21407 19125 21419 19128
rect 21361 19119 21419 19125
rect 22278 19116 22284 19128
rect 22336 19116 22342 19168
rect 552 19066 23368 19088
rect 552 19014 4322 19066
rect 4374 19014 4386 19066
rect 4438 19014 4450 19066
rect 4502 19014 4514 19066
rect 4566 19014 4578 19066
rect 4630 19014 23368 19066
rect 552 18992 23368 19014
rect 5994 18912 6000 18964
rect 6052 18912 6058 18964
rect 7009 18955 7067 18961
rect 7009 18921 7021 18955
rect 7055 18952 7067 18955
rect 7558 18952 7564 18964
rect 7055 18924 7564 18952
rect 7055 18921 7067 18924
rect 7009 18915 7067 18921
rect 7558 18912 7564 18924
rect 7616 18912 7622 18964
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 9125 18955 9183 18961
rect 8352 18924 8892 18952
rect 8352 18912 8358 18924
rect 6012 18884 6040 18912
rect 6457 18887 6515 18893
rect 5276 18856 6408 18884
rect 5276 18825 5304 18856
rect 5261 18819 5319 18825
rect 5261 18785 5273 18819
rect 5307 18785 5319 18819
rect 5261 18779 5319 18785
rect 5442 18776 5448 18828
rect 5500 18816 5506 18828
rect 5813 18819 5871 18825
rect 5813 18816 5825 18819
rect 5500 18788 5825 18816
rect 5500 18776 5506 18788
rect 5813 18785 5825 18788
rect 5859 18785 5871 18819
rect 5813 18779 5871 18785
rect 5997 18819 6055 18825
rect 5997 18785 6009 18819
rect 6043 18785 6055 18819
rect 5997 18779 6055 18785
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18748 5411 18751
rect 5534 18748 5540 18760
rect 5399 18720 5540 18748
rect 5399 18717 5411 18720
rect 5353 18711 5411 18717
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 5258 18640 5264 18692
rect 5316 18680 5322 18692
rect 6012 18680 6040 18779
rect 6270 18776 6276 18828
rect 6328 18776 6334 18828
rect 6380 18816 6408 18856
rect 6457 18853 6469 18887
rect 6503 18884 6515 18887
rect 8386 18884 8392 18896
rect 6503 18856 8392 18884
rect 6503 18853 6515 18856
rect 6457 18847 6515 18853
rect 6380 18788 6776 18816
rect 6638 18708 6644 18760
rect 6696 18708 6702 18760
rect 6748 18748 6776 18788
rect 6822 18776 6828 18828
rect 6880 18776 6886 18828
rect 7101 18819 7159 18825
rect 7101 18785 7113 18819
rect 7147 18816 7159 18819
rect 7190 18816 7196 18828
rect 7147 18788 7196 18816
rect 7147 18785 7159 18788
rect 7101 18779 7159 18785
rect 7190 18776 7196 18788
rect 7248 18776 7254 18828
rect 7300 18825 7328 18856
rect 8386 18844 8392 18856
rect 8444 18844 8450 18896
rect 8864 18828 8892 18924
rect 9125 18921 9137 18955
rect 9171 18952 9183 18955
rect 11238 18952 11244 18964
rect 9171 18924 11244 18952
rect 9171 18921 9183 18924
rect 9125 18915 9183 18921
rect 11238 18912 11244 18924
rect 11296 18912 11302 18964
rect 14277 18955 14335 18961
rect 14277 18921 14289 18955
rect 14323 18952 14335 18955
rect 14458 18952 14464 18964
rect 14323 18924 14464 18952
rect 14323 18921 14335 18924
rect 14277 18915 14335 18921
rect 14458 18912 14464 18924
rect 14516 18952 14522 18964
rect 14516 18924 15516 18952
rect 14516 18912 14522 18924
rect 10042 18844 10048 18896
rect 10100 18844 10106 18896
rect 12066 18844 12072 18896
rect 12124 18844 12130 18896
rect 13909 18887 13967 18893
rect 13909 18853 13921 18887
rect 13955 18853 13967 18887
rect 14642 18884 14648 18896
rect 13909 18847 13967 18853
rect 14476 18856 14648 18884
rect 7285 18819 7343 18825
rect 7285 18785 7297 18819
rect 7331 18785 7343 18819
rect 7285 18779 7343 18785
rect 7466 18776 7472 18828
rect 7524 18776 7530 18828
rect 8846 18776 8852 18828
rect 8904 18776 8910 18828
rect 8938 18776 8944 18828
rect 8996 18776 9002 18828
rect 9398 18776 9404 18828
rect 9456 18816 9462 18828
rect 9585 18819 9643 18825
rect 9585 18816 9597 18819
rect 9456 18788 9597 18816
rect 9456 18776 9462 18788
rect 9585 18785 9597 18788
rect 9631 18785 9643 18819
rect 9585 18779 9643 18785
rect 9861 18819 9919 18825
rect 9861 18785 9873 18819
rect 9907 18785 9919 18819
rect 9861 18779 9919 18785
rect 7742 18748 7748 18760
rect 6748 18720 7748 18748
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 8481 18751 8539 18757
rect 8481 18717 8493 18751
rect 8527 18748 8539 18751
rect 8754 18748 8760 18760
rect 8527 18720 8760 18748
rect 8527 18717 8539 18720
rect 8481 18711 8539 18717
rect 8754 18708 8760 18720
rect 8812 18708 8818 18760
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 9876 18748 9904 18779
rect 10594 18776 10600 18828
rect 10652 18776 10658 18828
rect 10962 18776 10968 18828
rect 11020 18776 11026 18828
rect 11330 18776 11336 18828
rect 11388 18776 11394 18828
rect 11698 18776 11704 18828
rect 11756 18816 11762 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11756 18788 11805 18816
rect 11756 18776 11762 18788
rect 11793 18785 11805 18788
rect 11839 18816 11851 18819
rect 12345 18819 12403 18825
rect 12345 18816 12357 18819
rect 11839 18788 12357 18816
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 12345 18785 12357 18788
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 13630 18776 13636 18828
rect 13688 18776 13694 18828
rect 13722 18776 13728 18828
rect 13780 18776 13786 18828
rect 13924 18816 13952 18847
rect 14185 18819 14243 18825
rect 14185 18816 14197 18819
rect 13924 18788 14197 18816
rect 14185 18785 14197 18788
rect 14231 18785 14243 18819
rect 14185 18779 14243 18785
rect 14366 18776 14372 18828
rect 14424 18816 14430 18828
rect 14476 18825 14504 18856
rect 14642 18844 14648 18856
rect 14700 18844 14706 18896
rect 14461 18819 14519 18825
rect 14461 18816 14473 18819
rect 14424 18788 14473 18816
rect 14424 18776 14430 18788
rect 14461 18785 14473 18788
rect 14507 18785 14519 18819
rect 14461 18779 14519 18785
rect 14734 18776 14740 18828
rect 14792 18776 14798 18828
rect 15102 18776 15108 18828
rect 15160 18816 15166 18828
rect 15197 18819 15255 18825
rect 15197 18816 15209 18819
rect 15160 18788 15209 18816
rect 15160 18776 15166 18788
rect 15197 18785 15209 18788
rect 15243 18816 15255 18819
rect 15378 18816 15384 18828
rect 15243 18788 15384 18816
rect 15243 18785 15255 18788
rect 15197 18779 15255 18785
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 15488 18825 15516 18924
rect 20530 18912 20536 18964
rect 20588 18952 20594 18964
rect 22370 18952 22376 18964
rect 20588 18924 22376 18952
rect 20588 18912 20594 18924
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 22554 18912 22560 18964
rect 22612 18952 22618 18964
rect 22649 18955 22707 18961
rect 22649 18952 22661 18955
rect 22612 18924 22661 18952
rect 22612 18912 22618 18924
rect 22649 18921 22661 18924
rect 22695 18921 22707 18955
rect 22649 18915 22707 18921
rect 16390 18844 16396 18896
rect 16448 18884 16454 18896
rect 16448 18856 16528 18884
rect 16448 18844 16454 18856
rect 16500 18825 16528 18856
rect 18230 18844 18236 18896
rect 18288 18884 18294 18896
rect 19788 18887 19846 18893
rect 18288 18856 18828 18884
rect 18288 18844 18294 18856
rect 15473 18819 15531 18825
rect 15473 18785 15485 18819
rect 15519 18785 15531 18819
rect 15473 18779 15531 18785
rect 16485 18819 16543 18825
rect 16485 18785 16497 18819
rect 16531 18785 16543 18819
rect 16485 18779 16543 18785
rect 18690 18776 18696 18828
rect 18748 18776 18754 18828
rect 18800 18825 18828 18856
rect 19788 18853 19800 18887
rect 19834 18884 19846 18887
rect 19978 18884 19984 18896
rect 19834 18856 19984 18884
rect 19834 18853 19846 18856
rect 19788 18847 19846 18853
rect 19978 18844 19984 18856
rect 20036 18844 20042 18896
rect 21266 18844 21272 18896
rect 21324 18884 21330 18896
rect 21514 18887 21572 18893
rect 21514 18884 21526 18887
rect 21324 18856 21526 18884
rect 21324 18844 21330 18856
rect 21514 18853 21526 18856
rect 21560 18853 21572 18887
rect 21514 18847 21572 18853
rect 18785 18819 18843 18825
rect 18785 18785 18797 18819
rect 18831 18785 18843 18819
rect 18785 18779 18843 18785
rect 18969 18819 19027 18825
rect 18969 18785 18981 18819
rect 19015 18785 19027 18819
rect 18969 18779 19027 18785
rect 9548 18720 9904 18748
rect 9548 18708 9554 18720
rect 10318 18708 10324 18760
rect 10376 18748 10382 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 10376 18720 10425 18748
rect 10376 18708 10382 18720
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 11974 18708 11980 18760
rect 12032 18748 12038 18760
rect 12253 18751 12311 18757
rect 12253 18748 12265 18751
rect 12032 18720 12265 18748
rect 12032 18708 12038 18720
rect 12253 18717 12265 18720
rect 12299 18717 12311 18751
rect 12253 18711 12311 18717
rect 13909 18751 13967 18757
rect 13909 18717 13921 18751
rect 13955 18717 13967 18751
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 13909 18711 13967 18717
rect 14384 18720 14657 18748
rect 5316 18652 6040 18680
rect 12713 18683 12771 18689
rect 5316 18640 5322 18652
rect 12713 18649 12725 18683
rect 12759 18680 12771 18683
rect 13814 18680 13820 18692
rect 12759 18652 13820 18680
rect 12759 18649 12771 18652
rect 12713 18643 12771 18649
rect 13814 18640 13820 18652
rect 13872 18680 13878 18692
rect 13924 18680 13952 18711
rect 13872 18652 13952 18680
rect 13872 18640 13878 18652
rect 5537 18615 5595 18621
rect 5537 18581 5549 18615
rect 5583 18612 5595 18615
rect 6730 18612 6736 18624
rect 5583 18584 6736 18612
rect 5583 18581 5595 18584
rect 5537 18575 5595 18581
rect 6730 18572 6736 18584
rect 6788 18572 6794 18624
rect 9309 18615 9367 18621
rect 9309 18581 9321 18615
rect 9355 18612 9367 18615
rect 9398 18612 9404 18624
rect 9355 18584 9404 18612
rect 9355 18581 9367 18584
rect 9309 18575 9367 18581
rect 9398 18572 9404 18584
rect 9456 18572 9462 18624
rect 10042 18572 10048 18624
rect 10100 18612 10106 18624
rect 10229 18615 10287 18621
rect 10229 18612 10241 18615
rect 10100 18584 10241 18612
rect 10100 18572 10106 18584
rect 10229 18581 10241 18584
rect 10275 18581 10287 18615
rect 10229 18575 10287 18581
rect 10781 18615 10839 18621
rect 10781 18581 10793 18615
rect 10827 18612 10839 18615
rect 11606 18612 11612 18624
rect 10827 18584 11612 18612
rect 10827 18581 10839 18584
rect 10781 18575 10839 18581
rect 11606 18572 11612 18584
rect 11664 18572 11670 18624
rect 14384 18612 14412 18720
rect 14645 18717 14657 18720
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 16298 18708 16304 18760
rect 16356 18748 16362 18760
rect 16393 18751 16451 18757
rect 16393 18748 16405 18751
rect 16356 18720 16405 18748
rect 16356 18708 16362 18720
rect 16393 18717 16405 18720
rect 16439 18717 16451 18751
rect 16393 18711 16451 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18748 18475 18751
rect 18506 18748 18512 18760
rect 18463 18720 18512 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 18506 18708 18512 18720
rect 18564 18708 18570 18760
rect 18708 18748 18736 18776
rect 18874 18748 18880 18760
rect 18708 18720 18880 18748
rect 18874 18708 18880 18720
rect 18932 18748 18938 18760
rect 18984 18748 19012 18779
rect 21910 18776 21916 18828
rect 21968 18816 21974 18828
rect 22833 18819 22891 18825
rect 22833 18816 22845 18819
rect 21968 18788 22845 18816
rect 21968 18776 21974 18788
rect 22833 18785 22845 18788
rect 22879 18785 22891 18819
rect 22833 18779 22891 18785
rect 22922 18776 22928 18828
rect 22980 18776 22986 18828
rect 18932 18720 19012 18748
rect 18932 18708 18938 18720
rect 19518 18708 19524 18760
rect 19576 18708 19582 18760
rect 21269 18751 21327 18757
rect 21269 18717 21281 18751
rect 21315 18717 21327 18751
rect 21269 18711 21327 18717
rect 14458 18640 14464 18692
rect 14516 18640 14522 18692
rect 15657 18683 15715 18689
rect 15657 18680 15669 18683
rect 14927 18652 15669 18680
rect 14927 18612 14955 18652
rect 15657 18649 15669 18652
rect 15703 18649 15715 18683
rect 15657 18643 15715 18649
rect 16114 18640 16120 18692
rect 16172 18640 16178 18692
rect 14384 18584 14955 18612
rect 15010 18572 15016 18624
rect 15068 18572 15074 18624
rect 15102 18572 15108 18624
rect 15160 18612 15166 18624
rect 15289 18615 15347 18621
rect 15289 18612 15301 18615
rect 15160 18584 15301 18612
rect 15160 18572 15166 18584
rect 15289 18581 15301 18584
rect 15335 18581 15347 18615
rect 15289 18575 15347 18581
rect 18506 18572 18512 18624
rect 18564 18572 18570 18624
rect 18601 18615 18659 18621
rect 18601 18581 18613 18615
rect 18647 18612 18659 18615
rect 18690 18612 18696 18624
rect 18647 18584 18696 18612
rect 18647 18581 18659 18584
rect 18601 18575 18659 18581
rect 18690 18572 18696 18584
rect 18748 18572 18754 18624
rect 18782 18572 18788 18624
rect 18840 18572 18846 18624
rect 20898 18572 20904 18624
rect 20956 18572 20962 18624
rect 21284 18612 21312 18711
rect 21542 18612 21548 18624
rect 21284 18584 21548 18612
rect 21542 18572 21548 18584
rect 21600 18572 21606 18624
rect 552 18522 23368 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 23368 18522
rect 552 18448 23368 18470
rect 4433 18411 4491 18417
rect 4433 18377 4445 18411
rect 4479 18408 4491 18411
rect 5626 18408 5632 18420
rect 4479 18380 5632 18408
rect 4479 18377 4491 18380
rect 4433 18371 4491 18377
rect 5626 18368 5632 18380
rect 5684 18368 5690 18420
rect 6822 18368 6828 18420
rect 6880 18408 6886 18420
rect 7929 18411 7987 18417
rect 7929 18408 7941 18411
rect 6880 18380 7941 18408
rect 6880 18368 6886 18380
rect 7929 18377 7941 18380
rect 7975 18377 7987 18411
rect 7929 18371 7987 18377
rect 8754 18368 8760 18420
rect 8812 18368 8818 18420
rect 10321 18411 10379 18417
rect 10321 18377 10333 18411
rect 10367 18408 10379 18411
rect 10410 18408 10416 18420
rect 10367 18380 10416 18408
rect 10367 18377 10379 18380
rect 10321 18371 10379 18377
rect 10410 18368 10416 18380
rect 10468 18408 10474 18420
rect 11330 18408 11336 18420
rect 10468 18380 11336 18408
rect 10468 18368 10474 18380
rect 11330 18368 11336 18380
rect 11388 18368 11394 18420
rect 11609 18411 11667 18417
rect 11609 18377 11621 18411
rect 11655 18408 11667 18411
rect 11655 18380 12434 18408
rect 11655 18377 11667 18380
rect 11609 18371 11667 18377
rect 6748 18312 7972 18340
rect 6748 18284 6776 18312
rect 5258 18232 5264 18284
rect 5316 18232 5322 18284
rect 6730 18232 6736 18284
rect 6788 18232 6794 18284
rect 7006 18272 7012 18284
rect 6840 18244 7012 18272
rect 4525 18207 4583 18213
rect 4525 18173 4537 18207
rect 4571 18204 4583 18207
rect 4571 18176 4660 18204
rect 4571 18173 4583 18176
rect 4525 18167 4583 18173
rect 4632 18145 4660 18176
rect 4798 18164 4804 18216
rect 4856 18204 4862 18216
rect 5169 18207 5227 18213
rect 5169 18204 5181 18207
rect 4856 18176 5181 18204
rect 4856 18164 4862 18176
rect 5169 18173 5181 18176
rect 5215 18204 5227 18207
rect 5442 18204 5448 18216
rect 5215 18176 5448 18204
rect 5215 18173 5227 18176
rect 5169 18167 5227 18173
rect 5442 18164 5448 18176
rect 5500 18164 5506 18216
rect 5905 18207 5963 18213
rect 5905 18173 5917 18207
rect 5951 18204 5963 18207
rect 5994 18204 6000 18216
rect 5951 18176 6000 18204
rect 5951 18173 5963 18176
rect 5905 18167 5963 18173
rect 5994 18164 6000 18176
rect 6052 18164 6058 18216
rect 6840 18213 6868 18244
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 7190 18232 7196 18284
rect 7248 18232 7254 18284
rect 7282 18232 7288 18284
rect 7340 18232 7346 18284
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7392 18244 7849 18272
rect 6181 18207 6239 18213
rect 6181 18173 6193 18207
rect 6227 18173 6239 18207
rect 6181 18167 6239 18173
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18173 6883 18207
rect 7392 18204 7420 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 6825 18167 6883 18173
rect 6932 18176 7420 18204
rect 7653 18207 7711 18213
rect 4617 18139 4675 18145
rect 4617 18105 4629 18139
rect 4663 18136 4675 18139
rect 4706 18136 4712 18148
rect 4663 18108 4712 18136
rect 4663 18105 4675 18108
rect 4617 18099 4675 18105
rect 4706 18096 4712 18108
rect 4764 18136 4770 18148
rect 5350 18136 5356 18148
rect 4764 18108 5356 18136
rect 4764 18096 4770 18108
rect 5350 18096 5356 18108
rect 5408 18096 5414 18148
rect 6196 18136 6224 18167
rect 6362 18136 6368 18148
rect 6196 18108 6368 18136
rect 6362 18096 6368 18108
rect 6420 18136 6426 18148
rect 6932 18136 6960 18176
rect 7653 18173 7665 18207
rect 7699 18204 7711 18207
rect 7742 18204 7748 18216
rect 7699 18176 7748 18204
rect 7699 18173 7711 18176
rect 7653 18167 7711 18173
rect 7742 18164 7748 18176
rect 7800 18164 7806 18216
rect 7944 18213 7972 18312
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8772 18272 8800 18368
rect 9493 18343 9551 18349
rect 9493 18309 9505 18343
rect 9539 18340 9551 18343
rect 10594 18340 10600 18352
rect 9539 18312 10600 18340
rect 9539 18309 9551 18312
rect 9493 18303 9551 18309
rect 10594 18300 10600 18312
rect 10652 18340 10658 18352
rect 10652 18312 10916 18340
rect 10652 18300 10658 18312
rect 10888 18281 10916 18312
rect 10962 18300 10968 18352
rect 11020 18340 11026 18352
rect 11698 18340 11704 18352
rect 11020 18312 11704 18340
rect 11020 18300 11026 18312
rect 11698 18300 11704 18312
rect 11756 18340 11762 18352
rect 12161 18343 12219 18349
rect 12161 18340 12173 18343
rect 11756 18312 12173 18340
rect 11756 18300 11762 18312
rect 12161 18309 12173 18312
rect 12207 18309 12219 18343
rect 12406 18340 12434 18380
rect 14550 18368 14556 18420
rect 14608 18408 14614 18420
rect 15197 18411 15255 18417
rect 15197 18408 15209 18411
rect 14608 18380 15209 18408
rect 14608 18368 14614 18380
rect 15197 18377 15209 18380
rect 15243 18377 15255 18411
rect 15197 18371 15255 18377
rect 18509 18411 18567 18417
rect 18509 18377 18521 18411
rect 18555 18408 18567 18411
rect 19794 18408 19800 18420
rect 18555 18380 19800 18408
rect 18555 18377 18567 18380
rect 18509 18371 18567 18377
rect 19794 18368 19800 18380
rect 19852 18368 19858 18420
rect 20349 18411 20407 18417
rect 20349 18377 20361 18411
rect 20395 18408 20407 18411
rect 20438 18408 20444 18420
rect 20395 18380 20444 18408
rect 20395 18377 20407 18380
rect 20349 18371 20407 18377
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 21085 18411 21143 18417
rect 21085 18377 21097 18411
rect 21131 18408 21143 18411
rect 21634 18408 21640 18420
rect 21131 18380 21640 18408
rect 21131 18377 21143 18380
rect 21085 18371 21143 18377
rect 21634 18368 21640 18380
rect 21692 18368 21698 18420
rect 13262 18340 13268 18352
rect 12406 18312 13268 18340
rect 12161 18303 12219 18309
rect 13262 18300 13268 18312
rect 13320 18300 13326 18352
rect 14366 18300 14372 18352
rect 14424 18340 14430 18352
rect 14424 18312 15240 18340
rect 14424 18300 14430 18312
rect 10873 18275 10931 18281
rect 8076 18244 8616 18272
rect 8772 18244 9260 18272
rect 8076 18232 8082 18244
rect 7929 18207 7987 18213
rect 7929 18173 7941 18207
rect 7975 18173 7987 18207
rect 7929 18167 7987 18173
rect 8110 18164 8116 18216
rect 8168 18164 8174 18216
rect 8386 18164 8392 18216
rect 8444 18164 8450 18216
rect 8588 18213 8616 18244
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18173 8631 18207
rect 8573 18167 8631 18173
rect 8846 18164 8852 18216
rect 8904 18204 8910 18216
rect 8941 18207 8999 18213
rect 8941 18204 8953 18207
rect 8904 18176 8953 18204
rect 8904 18164 8910 18176
rect 8941 18173 8953 18176
rect 8987 18173 8999 18207
rect 8941 18167 8999 18173
rect 6420 18108 6960 18136
rect 8956 18136 8984 18167
rect 9030 18164 9036 18216
rect 9088 18204 9094 18216
rect 9232 18213 9260 18244
rect 9324 18244 10272 18272
rect 9324 18213 9352 18244
rect 9125 18207 9183 18213
rect 9125 18204 9137 18207
rect 9088 18176 9137 18204
rect 9088 18164 9094 18176
rect 9125 18173 9137 18176
rect 9171 18173 9183 18207
rect 9125 18167 9183 18173
rect 9217 18207 9275 18213
rect 9217 18173 9229 18207
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 9309 18207 9367 18213
rect 9309 18173 9321 18207
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 9585 18207 9643 18213
rect 9585 18173 9597 18207
rect 9631 18173 9643 18207
rect 9585 18167 9643 18173
rect 9600 18136 9628 18167
rect 9766 18164 9772 18216
rect 9824 18164 9830 18216
rect 10244 18213 10272 18244
rect 10873 18241 10885 18275
rect 10919 18241 10931 18275
rect 10873 18235 10931 18241
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18272 11391 18275
rect 11793 18275 11851 18281
rect 11379 18244 11744 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 10229 18207 10287 18213
rect 10229 18173 10241 18207
rect 10275 18173 10287 18207
rect 10229 18167 10287 18173
rect 8956 18108 9628 18136
rect 10244 18136 10272 18167
rect 10318 18164 10324 18216
rect 10376 18204 10382 18216
rect 10965 18207 11023 18213
rect 10965 18204 10977 18207
rect 10376 18176 10977 18204
rect 10376 18164 10382 18176
rect 10965 18173 10977 18176
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 11606 18164 11612 18216
rect 11664 18164 11670 18216
rect 11716 18204 11744 18244
rect 11793 18241 11805 18275
rect 11839 18272 11851 18275
rect 14829 18275 14887 18281
rect 11839 18244 12388 18272
rect 11839 18241 11851 18244
rect 11793 18235 11851 18241
rect 12360 18216 12388 18244
rect 14829 18241 14841 18275
rect 14875 18272 14887 18275
rect 15010 18272 15016 18284
rect 14875 18244 15016 18272
rect 14875 18241 14887 18244
rect 14829 18235 14887 18241
rect 15010 18232 15016 18244
rect 15068 18232 15074 18284
rect 15105 18275 15163 18281
rect 15105 18241 15117 18275
rect 15151 18241 15163 18275
rect 15105 18235 15163 18241
rect 11974 18204 11980 18216
rect 11716 18176 11980 18204
rect 11974 18164 11980 18176
rect 12032 18164 12038 18216
rect 12069 18207 12127 18213
rect 12069 18173 12081 18207
rect 12115 18173 12127 18207
rect 12069 18167 12127 18173
rect 11054 18136 11060 18148
rect 10244 18108 11060 18136
rect 6420 18096 6426 18108
rect 11054 18096 11060 18108
rect 11112 18096 11118 18148
rect 11882 18096 11888 18148
rect 11940 18136 11946 18148
rect 12084 18136 12112 18167
rect 12342 18164 12348 18216
rect 12400 18164 12406 18216
rect 14737 18207 14795 18213
rect 14737 18173 14749 18207
rect 14783 18204 14795 18207
rect 14918 18204 14924 18216
rect 14783 18176 14924 18204
rect 14783 18173 14795 18176
rect 14737 18167 14795 18173
rect 14918 18164 14924 18176
rect 14976 18164 14982 18216
rect 15120 18204 15148 18235
rect 15212 18213 15240 18312
rect 18598 18300 18604 18352
rect 18656 18340 18662 18352
rect 19061 18343 19119 18349
rect 19061 18340 19073 18343
rect 18656 18312 19073 18340
rect 18656 18300 18662 18312
rect 19061 18309 19073 18312
rect 19107 18309 19119 18343
rect 19061 18303 19119 18309
rect 21545 18343 21603 18349
rect 21545 18309 21557 18343
rect 21591 18309 21603 18343
rect 21545 18303 21603 18309
rect 15746 18232 15752 18284
rect 15804 18272 15810 18284
rect 16209 18275 16267 18281
rect 16209 18272 16221 18275
rect 15804 18244 16221 18272
rect 15804 18232 15810 18244
rect 16209 18241 16221 18244
rect 16255 18272 16267 18275
rect 18616 18272 18644 18300
rect 16255 18244 16988 18272
rect 16255 18241 16267 18244
rect 16209 18235 16267 18241
rect 15028 18176 15148 18204
rect 15197 18207 15255 18213
rect 11940 18108 12112 18136
rect 15028 18136 15056 18176
rect 15197 18173 15209 18207
rect 15243 18173 15255 18207
rect 15197 18167 15255 18173
rect 15378 18164 15384 18216
rect 15436 18164 15442 18216
rect 15654 18164 15660 18216
rect 15712 18204 15718 18216
rect 16114 18204 16120 18216
rect 15712 18176 16120 18204
rect 15712 18164 15718 18176
rect 16114 18164 16120 18176
rect 16172 18204 16178 18216
rect 16960 18213 16988 18244
rect 18156 18244 18644 18272
rect 16301 18207 16359 18213
rect 16301 18204 16313 18207
rect 16172 18176 16313 18204
rect 16172 18164 16178 18176
rect 16301 18173 16313 18176
rect 16347 18204 16359 18207
rect 16761 18207 16819 18213
rect 16761 18204 16773 18207
rect 16347 18176 16773 18204
rect 16347 18173 16359 18176
rect 16301 18167 16359 18173
rect 16761 18173 16773 18176
rect 16807 18173 16819 18207
rect 16761 18167 16819 18173
rect 16945 18207 17003 18213
rect 16945 18173 16957 18207
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 17494 18164 17500 18216
rect 17552 18164 17558 18216
rect 17678 18164 17684 18216
rect 17736 18164 17742 18216
rect 18156 18213 18184 18244
rect 18690 18232 18696 18284
rect 18748 18272 18754 18284
rect 18966 18272 18972 18284
rect 18748 18244 18972 18272
rect 18748 18232 18754 18244
rect 18966 18232 18972 18244
rect 19024 18232 19030 18284
rect 20717 18275 20775 18281
rect 20717 18241 20729 18275
rect 20763 18272 20775 18275
rect 20898 18272 20904 18284
rect 20763 18244 20904 18272
rect 20763 18241 20775 18244
rect 20717 18235 20775 18241
rect 20898 18232 20904 18244
rect 20956 18232 20962 18284
rect 21560 18272 21588 18303
rect 21560 18244 21772 18272
rect 17865 18207 17923 18213
rect 17865 18173 17877 18207
rect 17911 18173 17923 18207
rect 17865 18167 17923 18173
rect 18141 18207 18199 18213
rect 18141 18173 18153 18207
rect 18187 18173 18199 18207
rect 18141 18167 18199 18173
rect 18509 18207 18567 18213
rect 18509 18173 18521 18207
rect 18555 18204 18567 18207
rect 18598 18204 18604 18216
rect 18555 18176 18604 18204
rect 18555 18173 18567 18176
rect 18509 18167 18567 18173
rect 15470 18136 15476 18148
rect 15028 18108 15476 18136
rect 11940 18096 11946 18108
rect 15470 18096 15476 18108
rect 15528 18096 15534 18148
rect 17586 18096 17592 18148
rect 17644 18136 17650 18148
rect 17880 18136 17908 18167
rect 18598 18164 18604 18176
rect 18656 18204 18662 18216
rect 18782 18204 18788 18216
rect 18656 18176 18788 18204
rect 18656 18164 18662 18176
rect 18782 18164 18788 18176
rect 18840 18164 18846 18216
rect 18874 18164 18880 18216
rect 18932 18164 18938 18216
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18204 19211 18207
rect 19334 18204 19340 18216
rect 19199 18176 19340 18204
rect 19199 18173 19211 18176
rect 19153 18167 19211 18173
rect 19334 18164 19340 18176
rect 19392 18164 19398 18216
rect 20530 18164 20536 18216
rect 20588 18204 20594 18216
rect 20993 18207 21051 18213
rect 20993 18204 21005 18207
rect 20588 18176 21005 18204
rect 20588 18164 20594 18176
rect 20993 18173 21005 18176
rect 21039 18173 21051 18207
rect 20993 18167 21051 18173
rect 21266 18164 21272 18216
rect 21324 18164 21330 18216
rect 21634 18164 21640 18216
rect 21692 18164 21698 18216
rect 21744 18204 21772 18244
rect 21893 18207 21951 18213
rect 21893 18204 21905 18207
rect 21744 18176 21905 18204
rect 21893 18173 21905 18176
rect 21939 18173 21951 18207
rect 21893 18167 21951 18173
rect 17644 18108 17908 18136
rect 17644 18096 17650 18108
rect 21542 18096 21548 18148
rect 21600 18096 21606 18148
rect 5169 18071 5227 18077
rect 5169 18037 5181 18071
rect 5215 18068 5227 18071
rect 6270 18068 6276 18080
rect 5215 18040 6276 18068
rect 5215 18037 5227 18040
rect 5169 18031 5227 18037
rect 6270 18028 6276 18040
rect 6328 18028 6334 18080
rect 6546 18028 6552 18080
rect 6604 18028 6610 18080
rect 7098 18028 7104 18080
rect 7156 18068 7162 18080
rect 7377 18071 7435 18077
rect 7377 18068 7389 18071
rect 7156 18040 7389 18068
rect 7156 18028 7162 18040
rect 7377 18037 7389 18040
rect 7423 18068 7435 18071
rect 8110 18068 8116 18080
rect 7423 18040 8116 18068
rect 7423 18037 7435 18040
rect 7377 18031 7435 18037
rect 8110 18028 8116 18040
rect 8168 18028 8174 18080
rect 9769 18071 9827 18077
rect 9769 18037 9781 18071
rect 9815 18068 9827 18071
rect 9858 18068 9864 18080
rect 9815 18040 9864 18068
rect 9815 18037 9827 18040
rect 9769 18031 9827 18037
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 15562 18028 15568 18080
rect 15620 18028 15626 18080
rect 16669 18071 16727 18077
rect 16669 18037 16681 18071
rect 16715 18068 16727 18071
rect 16758 18068 16764 18080
rect 16715 18040 16764 18068
rect 16715 18037 16727 18040
rect 16669 18031 16727 18037
rect 16758 18028 16764 18040
rect 16816 18028 16822 18080
rect 16850 18028 16856 18080
rect 16908 18028 16914 18080
rect 18690 18028 18696 18080
rect 18748 18028 18754 18080
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 21910 18068 21916 18080
rect 21407 18040 21916 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 22370 18028 22376 18080
rect 22428 18068 22434 18080
rect 22922 18068 22928 18080
rect 22428 18040 22928 18068
rect 22428 18028 22434 18040
rect 22922 18028 22928 18040
rect 22980 18068 22986 18080
rect 23017 18071 23075 18077
rect 23017 18068 23029 18071
rect 22980 18040 23029 18068
rect 22980 18028 22986 18040
rect 23017 18037 23029 18040
rect 23063 18037 23075 18071
rect 23017 18031 23075 18037
rect 552 17978 23368 18000
rect 552 17926 4322 17978
rect 4374 17926 4386 17978
rect 4438 17926 4450 17978
rect 4502 17926 4514 17978
rect 4566 17926 4578 17978
rect 4630 17926 23368 17978
rect 552 17904 23368 17926
rect 5166 17864 5172 17876
rect 4632 17836 5172 17864
rect 4632 17805 4660 17836
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 5629 17867 5687 17873
rect 5629 17864 5641 17867
rect 5592 17836 5641 17864
rect 5592 17824 5598 17836
rect 5629 17833 5641 17836
rect 5675 17833 5687 17867
rect 5629 17827 5687 17833
rect 8665 17867 8723 17873
rect 8665 17833 8677 17867
rect 8711 17833 8723 17867
rect 8665 17827 8723 17833
rect 4617 17799 4675 17805
rect 4617 17765 4629 17799
rect 4663 17765 4675 17799
rect 4617 17759 4675 17765
rect 4798 17756 4804 17808
rect 4856 17756 4862 17808
rect 4985 17799 5043 17805
rect 4985 17765 4997 17799
rect 5031 17796 5043 17799
rect 5258 17796 5264 17808
rect 5031 17768 5264 17796
rect 5031 17765 5043 17768
rect 4985 17759 5043 17765
rect 5258 17756 5264 17768
rect 5316 17796 5322 17808
rect 5813 17799 5871 17805
rect 5813 17796 5825 17799
rect 5316 17768 5825 17796
rect 5316 17756 5322 17768
rect 5813 17765 5825 17768
rect 5859 17765 5871 17799
rect 5813 17759 5871 17765
rect 7653 17799 7711 17805
rect 7653 17765 7665 17799
rect 7699 17796 7711 17799
rect 8680 17796 8708 17827
rect 10318 17824 10324 17876
rect 10376 17824 10382 17876
rect 13081 17867 13139 17873
rect 13081 17833 13093 17867
rect 13127 17833 13139 17867
rect 13081 17827 13139 17833
rect 10778 17796 10784 17808
rect 7699 17768 8616 17796
rect 8680 17768 10784 17796
rect 7699 17765 7711 17768
rect 7653 17759 7711 17765
rect 5077 17731 5135 17737
rect 5077 17697 5089 17731
rect 5123 17697 5135 17731
rect 5077 17691 5135 17697
rect 5092 17660 5120 17691
rect 5350 17688 5356 17740
rect 5408 17688 5414 17740
rect 5445 17731 5503 17737
rect 5445 17697 5457 17731
rect 5491 17728 5503 17731
rect 5626 17728 5632 17740
rect 5491 17700 5632 17728
rect 5491 17697 5503 17700
rect 5445 17691 5503 17697
rect 5626 17688 5632 17700
rect 5684 17688 5690 17740
rect 6181 17731 6239 17737
rect 6181 17728 6193 17731
rect 5736 17700 6193 17728
rect 5534 17660 5540 17672
rect 5092 17632 5540 17660
rect 5534 17620 5540 17632
rect 5592 17660 5598 17672
rect 5736 17660 5764 17700
rect 6181 17697 6193 17700
rect 6227 17728 6239 17731
rect 6270 17728 6276 17740
rect 6227 17700 6276 17728
rect 6227 17697 6239 17700
rect 6181 17691 6239 17697
rect 6270 17688 6276 17700
rect 6328 17688 6334 17740
rect 6546 17688 6552 17740
rect 6604 17728 6610 17740
rect 6825 17731 6883 17737
rect 6825 17728 6837 17731
rect 6604 17700 6837 17728
rect 6604 17688 6610 17700
rect 6825 17697 6837 17700
rect 6871 17697 6883 17731
rect 6825 17691 6883 17697
rect 8297 17731 8355 17737
rect 8297 17697 8309 17731
rect 8343 17728 8355 17731
rect 8588 17728 8616 17768
rect 10778 17756 10784 17768
rect 10836 17796 10842 17808
rect 13096 17796 13124 17827
rect 14458 17824 14464 17876
rect 14516 17864 14522 17876
rect 16022 17864 16028 17876
rect 14516 17836 16028 17864
rect 14516 17824 14522 17836
rect 16022 17824 16028 17836
rect 16080 17824 16086 17876
rect 16485 17867 16543 17873
rect 16485 17833 16497 17867
rect 16531 17864 16543 17867
rect 17678 17864 17684 17876
rect 16531 17836 17684 17864
rect 16531 17833 16543 17836
rect 16485 17827 16543 17833
rect 17678 17824 17684 17836
rect 17736 17824 17742 17876
rect 18141 17867 18199 17873
rect 18141 17833 18153 17867
rect 18187 17864 18199 17867
rect 18187 17836 18644 17864
rect 18187 17833 18199 17836
rect 18141 17827 18199 17833
rect 14001 17799 14059 17805
rect 14001 17796 14013 17799
rect 10836 17768 11192 17796
rect 13096 17768 14013 17796
rect 10836 17756 10842 17768
rect 9674 17728 9680 17740
rect 8343 17700 8524 17728
rect 8588 17700 9680 17728
rect 8343 17697 8355 17700
rect 8297 17691 8355 17697
rect 5592 17632 5764 17660
rect 5592 17620 5598 17632
rect 5994 17620 6000 17672
rect 6052 17620 6058 17672
rect 6733 17663 6791 17669
rect 6733 17660 6745 17663
rect 6196 17632 6745 17660
rect 6196 17601 6224 17632
rect 6733 17629 6745 17632
rect 6779 17660 6791 17663
rect 7006 17660 7012 17672
rect 6779 17632 7012 17660
rect 6779 17629 6791 17632
rect 6733 17623 6791 17629
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 7190 17620 7196 17672
rect 7248 17660 7254 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7248 17632 8217 17660
rect 7248 17620 7254 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8496 17660 8524 17700
rect 9674 17688 9680 17700
rect 9732 17728 9738 17740
rect 9953 17731 10011 17737
rect 9953 17728 9965 17731
rect 9732 17700 9965 17728
rect 9732 17688 9738 17700
rect 9953 17697 9965 17700
rect 9999 17728 10011 17731
rect 10226 17728 10232 17740
rect 9999 17700 10232 17728
rect 9999 17697 10011 17700
rect 9953 17691 10011 17697
rect 10226 17688 10232 17700
rect 10284 17688 10290 17740
rect 10962 17688 10968 17740
rect 11020 17688 11026 17740
rect 11164 17737 11192 17768
rect 11149 17731 11207 17737
rect 11149 17697 11161 17731
rect 11195 17697 11207 17731
rect 11149 17691 11207 17697
rect 12066 17688 12072 17740
rect 12124 17728 12130 17740
rect 12253 17731 12311 17737
rect 12253 17728 12265 17731
rect 12124 17700 12265 17728
rect 12124 17688 12130 17700
rect 12253 17697 12265 17700
rect 12299 17728 12311 17731
rect 12526 17728 12532 17740
rect 12299 17700 12532 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 12526 17688 12532 17700
rect 12584 17728 12590 17740
rect 13372 17737 13400 17768
rect 14001 17765 14013 17768
rect 14047 17765 14059 17799
rect 16114 17796 16120 17808
rect 14001 17759 14059 17765
rect 15856 17768 16120 17796
rect 12713 17731 12771 17737
rect 12713 17728 12725 17731
rect 12584 17700 12725 17728
rect 12584 17688 12590 17700
rect 12713 17697 12725 17700
rect 12759 17697 12771 17731
rect 12713 17691 12771 17697
rect 13357 17731 13415 17737
rect 13357 17697 13369 17731
rect 13403 17697 13415 17731
rect 13357 17691 13415 17697
rect 13817 17731 13875 17737
rect 13817 17697 13829 17731
rect 13863 17697 13875 17731
rect 13817 17691 13875 17697
rect 8570 17660 8576 17672
rect 8496 17632 8576 17660
rect 8205 17623 8263 17629
rect 8570 17620 8576 17632
rect 8628 17620 8634 17672
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 10134 17660 10140 17672
rect 10091 17632 10140 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17660 11115 17663
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 11103 17632 11713 17660
rect 11103 17629 11115 17632
rect 11057 17623 11115 17629
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11701 17623 11759 17629
rect 12342 17620 12348 17672
rect 12400 17660 12406 17672
rect 12621 17663 12679 17669
rect 12621 17660 12633 17663
rect 12400 17632 12633 17660
rect 12400 17620 12406 17632
rect 12621 17629 12633 17632
rect 12667 17629 12679 17663
rect 12621 17623 12679 17629
rect 13262 17620 13268 17672
rect 13320 17660 13326 17672
rect 13832 17660 13860 17691
rect 15654 17688 15660 17740
rect 15712 17688 15718 17740
rect 15746 17688 15752 17740
rect 15804 17688 15810 17740
rect 15764 17660 15792 17688
rect 13320 17632 13860 17660
rect 13924 17632 15792 17660
rect 13320 17620 13326 17632
rect 6181 17595 6239 17601
rect 6181 17561 6193 17595
rect 6227 17561 6239 17595
rect 6181 17555 6239 17561
rect 11977 17595 12035 17601
rect 11977 17561 11989 17595
rect 12023 17592 12035 17595
rect 13924 17592 13952 17632
rect 15856 17592 15884 17768
rect 16114 17756 16120 17768
rect 16172 17756 16178 17808
rect 16333 17799 16391 17805
rect 16333 17765 16345 17799
rect 16379 17796 16391 17799
rect 17126 17796 17132 17808
rect 16379 17768 17132 17796
rect 16379 17765 16391 17768
rect 16333 17759 16391 17765
rect 17126 17756 17132 17768
rect 17184 17756 17190 17808
rect 17604 17768 18368 17796
rect 15933 17731 15991 17737
rect 15933 17697 15945 17731
rect 15979 17728 15991 17731
rect 16761 17731 16819 17737
rect 16761 17728 16773 17731
rect 15979 17700 16773 17728
rect 15979 17697 15991 17700
rect 15933 17691 15991 17697
rect 16316 17672 16344 17700
rect 16761 17697 16773 17700
rect 16807 17697 16819 17731
rect 16761 17691 16819 17697
rect 16850 17688 16856 17740
rect 16908 17728 16914 17740
rect 17037 17731 17095 17737
rect 17037 17728 17049 17731
rect 16908 17700 17049 17728
rect 16908 17688 16914 17700
rect 17037 17697 17049 17700
rect 17083 17697 17095 17731
rect 17037 17691 17095 17697
rect 17221 17731 17279 17737
rect 17221 17697 17233 17731
rect 17267 17728 17279 17731
rect 17402 17728 17408 17740
rect 17267 17700 17408 17728
rect 17267 17697 17279 17700
rect 17221 17691 17279 17697
rect 17402 17688 17408 17700
rect 17460 17688 17466 17740
rect 17604 17737 17632 17768
rect 17589 17731 17647 17737
rect 17589 17697 17601 17731
rect 17635 17697 17647 17731
rect 17589 17691 17647 17697
rect 18049 17731 18107 17737
rect 18049 17697 18061 17731
rect 18095 17728 18107 17731
rect 18230 17728 18236 17740
rect 18095 17700 18236 17728
rect 18095 17697 18107 17700
rect 18049 17691 18107 17697
rect 16298 17620 16304 17672
rect 16356 17620 16362 17672
rect 16482 17620 16488 17672
rect 16540 17660 16546 17672
rect 16868 17660 16896 17688
rect 16540 17632 16896 17660
rect 16540 17620 16546 17632
rect 17310 17620 17316 17672
rect 17368 17660 17374 17672
rect 17604 17660 17632 17691
rect 18230 17688 18236 17700
rect 18288 17688 18294 17740
rect 18340 17737 18368 17768
rect 18506 17756 18512 17808
rect 18564 17756 18570 17808
rect 18616 17796 18644 17836
rect 21542 17824 21548 17876
rect 21600 17864 21606 17876
rect 21637 17867 21695 17873
rect 21637 17864 21649 17867
rect 21600 17836 21649 17864
rect 21600 17824 21606 17836
rect 21637 17833 21649 17836
rect 21683 17833 21695 17867
rect 21637 17827 21695 17833
rect 19030 17799 19088 17805
rect 19030 17796 19042 17799
rect 18616 17768 19042 17796
rect 19030 17765 19042 17768
rect 19076 17765 19088 17799
rect 19030 17759 19088 17765
rect 23014 17756 23020 17808
rect 23072 17756 23078 17808
rect 18325 17731 18383 17737
rect 18325 17697 18337 17731
rect 18371 17697 18383 17731
rect 18325 17691 18383 17697
rect 18417 17731 18475 17737
rect 18417 17697 18429 17731
rect 18463 17697 18475 17731
rect 18417 17691 18475 17697
rect 17368 17632 17632 17660
rect 17727 17663 17785 17669
rect 17368 17620 17374 17632
rect 17727 17629 17739 17663
rect 17773 17660 17785 17663
rect 18138 17660 18144 17672
rect 17773 17632 18144 17660
rect 17773 17629 17785 17632
rect 17727 17623 17785 17629
rect 18138 17620 18144 17632
rect 18196 17620 18202 17672
rect 12023 17564 13952 17592
rect 14108 17564 15884 17592
rect 12023 17561 12035 17564
rect 11977 17555 12035 17561
rect 5442 17484 5448 17536
rect 5500 17524 5506 17536
rect 6454 17524 6460 17536
rect 5500 17496 6460 17524
rect 5500 17484 5506 17496
rect 6454 17484 6460 17496
rect 6512 17484 6518 17536
rect 8846 17484 8852 17536
rect 8904 17524 8910 17536
rect 10042 17524 10048 17536
rect 8904 17496 10048 17524
rect 8904 17484 8910 17496
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 13725 17527 13783 17533
rect 13725 17493 13737 17527
rect 13771 17524 13783 17527
rect 14108 17524 14136 17564
rect 16022 17552 16028 17604
rect 16080 17592 16086 17604
rect 16577 17595 16635 17601
rect 16080 17564 16344 17592
rect 16080 17552 16086 17564
rect 13771 17496 14136 17524
rect 14185 17527 14243 17533
rect 13771 17493 13783 17496
rect 13725 17487 13783 17493
rect 14185 17493 14197 17527
rect 14231 17524 14243 17527
rect 16206 17524 16212 17536
rect 14231 17496 16212 17524
rect 14231 17493 14243 17496
rect 14185 17487 14243 17493
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 16316 17533 16344 17564
rect 16577 17561 16589 17595
rect 16623 17592 16635 17595
rect 17586 17592 17592 17604
rect 16623 17564 17592 17592
rect 16623 17561 16635 17564
rect 16577 17555 16635 17561
rect 17586 17552 17592 17564
rect 17644 17552 17650 17604
rect 17865 17595 17923 17601
rect 17865 17561 17877 17595
rect 17911 17592 17923 17595
rect 18322 17592 18328 17604
rect 17911 17564 18328 17592
rect 17911 17561 17923 17564
rect 17865 17555 17923 17561
rect 18322 17552 18328 17564
rect 18380 17552 18386 17604
rect 16301 17527 16359 17533
rect 16301 17493 16313 17527
rect 16347 17493 16359 17527
rect 16301 17487 16359 17493
rect 17957 17527 18015 17533
rect 17957 17493 17969 17527
rect 18003 17524 18015 17527
rect 18046 17524 18052 17536
rect 18003 17496 18052 17524
rect 18003 17493 18015 17496
rect 17957 17487 18015 17493
rect 18046 17484 18052 17496
rect 18104 17484 18110 17536
rect 18432 17524 18460 17691
rect 18690 17688 18696 17740
rect 18748 17688 18754 17740
rect 19518 17728 19524 17740
rect 18800 17700 19524 17728
rect 18800 17669 18828 17700
rect 19518 17688 19524 17700
rect 19576 17688 19582 17740
rect 21266 17688 21272 17740
rect 21324 17728 21330 17740
rect 21818 17728 21824 17740
rect 21324 17700 21824 17728
rect 21324 17688 21330 17700
rect 21818 17688 21824 17700
rect 21876 17688 21882 17740
rect 21910 17688 21916 17740
rect 21968 17688 21974 17740
rect 22370 17688 22376 17740
rect 22428 17688 22434 17740
rect 22554 17688 22560 17740
rect 22612 17688 22618 17740
rect 18785 17663 18843 17669
rect 18785 17660 18797 17663
rect 18708 17632 18797 17660
rect 18708 17604 18736 17632
rect 18785 17629 18797 17632
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 20806 17620 20812 17672
rect 20864 17660 20870 17672
rect 21637 17663 21695 17669
rect 21637 17660 21649 17663
rect 20864 17632 21649 17660
rect 20864 17620 20870 17632
rect 21637 17629 21649 17632
rect 21683 17660 21695 17663
rect 22186 17660 22192 17672
rect 21683 17632 22192 17660
rect 21683 17629 21695 17632
rect 21637 17623 21695 17629
rect 22186 17620 22192 17632
rect 22244 17620 22250 17672
rect 22281 17663 22339 17669
rect 22281 17629 22293 17663
rect 22327 17660 22339 17663
rect 22830 17660 22836 17672
rect 22327 17632 22836 17660
rect 22327 17629 22339 17632
rect 22281 17623 22339 17629
rect 18690 17552 18696 17604
rect 18748 17552 18754 17604
rect 22094 17552 22100 17604
rect 22152 17592 22158 17604
rect 22296 17592 22324 17623
rect 22830 17620 22836 17632
rect 22888 17620 22894 17672
rect 22152 17564 22324 17592
rect 22152 17552 22158 17564
rect 19426 17524 19432 17536
rect 18432 17496 19432 17524
rect 19426 17484 19432 17496
rect 19484 17524 19490 17536
rect 20165 17527 20223 17533
rect 20165 17524 20177 17527
rect 19484 17496 20177 17524
rect 19484 17484 19490 17496
rect 20165 17493 20177 17496
rect 20211 17493 20223 17527
rect 20165 17487 20223 17493
rect 552 17434 23368 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 23368 17434
rect 552 17360 23368 17382
rect 5994 17320 6000 17332
rect 5644 17292 6000 17320
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17184 5135 17187
rect 5123 17156 5488 17184
rect 5123 17153 5135 17156
rect 5077 17147 5135 17153
rect 5460 17128 5488 17156
rect 4890 17076 4896 17128
rect 4948 17076 4954 17128
rect 5258 17076 5264 17128
rect 5316 17076 5322 17128
rect 5350 17076 5356 17128
rect 5408 17076 5414 17128
rect 5442 17076 5448 17128
rect 5500 17076 5506 17128
rect 5644 17125 5672 17292
rect 5994 17280 6000 17292
rect 6052 17280 6058 17332
rect 6273 17323 6331 17329
rect 6273 17289 6285 17323
rect 6319 17320 6331 17323
rect 6914 17320 6920 17332
rect 6319 17292 6920 17320
rect 6319 17289 6331 17292
rect 6273 17283 6331 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 9490 17280 9496 17332
rect 9548 17320 9554 17332
rect 10962 17320 10968 17332
rect 9548 17292 10968 17320
rect 9548 17280 9554 17292
rect 5902 17212 5908 17264
rect 5960 17252 5966 17264
rect 6362 17252 6368 17264
rect 5960 17224 6368 17252
rect 5960 17212 5966 17224
rect 6362 17212 6368 17224
rect 6420 17212 6426 17264
rect 6549 17255 6607 17261
rect 6549 17221 6561 17255
rect 6595 17221 6607 17255
rect 6549 17215 6607 17221
rect 6564 17184 6592 17215
rect 9030 17212 9036 17264
rect 9088 17252 9094 17264
rect 9217 17255 9275 17261
rect 9217 17252 9229 17255
rect 9088 17224 9229 17252
rect 9088 17212 9094 17224
rect 9217 17221 9229 17224
rect 9263 17221 9275 17255
rect 9858 17252 9864 17264
rect 9217 17215 9275 17221
rect 9784 17224 9864 17252
rect 9784 17184 9812 17224
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 9968 17224 10364 17252
rect 9968 17184 9996 17224
rect 5736 17156 6592 17184
rect 8956 17156 9812 17184
rect 9888 17156 9996 17184
rect 5736 17125 5764 17156
rect 5603 17119 5672 17125
rect 5603 17085 5615 17119
rect 5649 17088 5672 17119
rect 5721 17119 5779 17125
rect 5649 17085 5661 17088
rect 5603 17079 5661 17085
rect 5721 17085 5733 17119
rect 5767 17085 5779 17119
rect 5721 17079 5779 17085
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17085 5963 17119
rect 6181 17119 6239 17125
rect 6181 17116 6193 17119
rect 5905 17079 5963 17085
rect 6104 17088 6193 17116
rect 5810 17008 5816 17060
rect 5868 17008 5874 17060
rect 5166 16940 5172 16992
rect 5224 16980 5230 16992
rect 5920 16980 5948 17079
rect 6104 16992 6132 17088
rect 6181 17085 6193 17088
rect 6227 17085 6239 17119
rect 6181 17079 6239 17085
rect 6362 17076 6368 17128
rect 6420 17076 6426 17128
rect 6454 17076 6460 17128
rect 6512 17076 6518 17128
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6604 17088 6837 17116
rect 6604 17076 6610 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7006 17076 7012 17128
rect 7064 17076 7070 17128
rect 8846 17076 8852 17128
rect 8904 17076 8910 17128
rect 8956 17125 8984 17156
rect 8941 17119 8999 17125
rect 8941 17085 8953 17119
rect 8987 17085 8999 17119
rect 9306 17116 9312 17128
rect 8941 17079 8999 17085
rect 9048 17088 9312 17116
rect 6917 17051 6975 17057
rect 6917 17017 6929 17051
rect 6963 17048 6975 17051
rect 9048 17048 9076 17088
rect 9306 17076 9312 17088
rect 9364 17116 9370 17128
rect 9401 17119 9459 17125
rect 9401 17116 9413 17119
rect 9364 17088 9413 17116
rect 9364 17076 9370 17088
rect 9401 17085 9413 17088
rect 9447 17085 9459 17119
rect 9401 17079 9459 17085
rect 9674 17076 9680 17128
rect 9732 17076 9738 17128
rect 9888 17125 9916 17156
rect 10226 17144 10232 17196
rect 10284 17144 10290 17196
rect 10336 17125 10364 17224
rect 10520 17184 10548 17292
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 11149 17323 11207 17329
rect 11149 17289 11161 17323
rect 11195 17320 11207 17323
rect 12342 17320 12348 17332
rect 11195 17292 12348 17320
rect 11195 17289 11207 17292
rect 11149 17283 11207 17289
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 15010 17280 15016 17332
rect 15068 17280 15074 17332
rect 16393 17323 16451 17329
rect 16393 17289 16405 17323
rect 16439 17289 16451 17323
rect 16393 17283 16451 17289
rect 14553 17255 14611 17261
rect 14553 17221 14565 17255
rect 14599 17252 14611 17255
rect 15378 17252 15384 17264
rect 14599 17224 15384 17252
rect 14599 17221 14611 17224
rect 14553 17215 14611 17221
rect 15378 17212 15384 17224
rect 15436 17212 15442 17264
rect 15473 17255 15531 17261
rect 15473 17221 15485 17255
rect 15519 17252 15531 17255
rect 16025 17255 16083 17261
rect 16025 17252 16037 17255
rect 15519 17224 16037 17252
rect 15519 17221 15531 17224
rect 15473 17215 15531 17221
rect 16025 17221 16037 17224
rect 16071 17221 16083 17255
rect 16408 17252 16436 17283
rect 17126 17280 17132 17332
rect 17184 17280 17190 17332
rect 17402 17280 17408 17332
rect 17460 17280 17466 17332
rect 17678 17280 17684 17332
rect 17736 17280 17742 17332
rect 18138 17280 18144 17332
rect 18196 17320 18202 17332
rect 18966 17320 18972 17332
rect 18196 17292 18972 17320
rect 18196 17280 18202 17292
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 22094 17320 22100 17332
rect 20824 17292 22100 17320
rect 16482 17252 16488 17264
rect 16408 17224 16488 17252
rect 16025 17215 16083 17221
rect 16482 17212 16488 17224
rect 16540 17212 16546 17264
rect 16942 17212 16948 17264
rect 17000 17212 17006 17264
rect 17957 17255 18015 17261
rect 17957 17221 17969 17255
rect 18003 17221 18015 17255
rect 17957 17215 18015 17221
rect 10689 17187 10747 17193
rect 10689 17184 10701 17187
rect 10520 17156 10701 17184
rect 10689 17153 10701 17156
rect 10735 17153 10747 17187
rect 15562 17184 15568 17196
rect 10689 17147 10747 17153
rect 14568 17156 15568 17184
rect 9861 17119 9919 17125
rect 9861 17085 9873 17119
rect 9907 17085 9919 17119
rect 9861 17079 9919 17085
rect 10321 17119 10379 17125
rect 10321 17085 10333 17119
rect 10367 17116 10379 17119
rect 10410 17116 10416 17128
rect 10367 17088 10416 17116
rect 10367 17085 10379 17088
rect 10321 17079 10379 17085
rect 10410 17076 10416 17088
rect 10468 17076 10474 17128
rect 10778 17076 10784 17128
rect 10836 17076 10842 17128
rect 14568 17125 14596 17156
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 16298 17144 16304 17196
rect 16356 17144 16362 17196
rect 16850 17144 16856 17196
rect 16908 17184 16914 17196
rect 17494 17184 17500 17196
rect 16908 17156 17500 17184
rect 16908 17144 16914 17156
rect 17494 17144 17500 17156
rect 17552 17184 17558 17196
rect 17681 17187 17739 17193
rect 17681 17184 17693 17187
rect 17552 17156 17693 17184
rect 17552 17144 17558 17156
rect 17681 17153 17693 17156
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 14277 17119 14335 17125
rect 14277 17085 14289 17119
rect 14323 17085 14335 17119
rect 14277 17079 14335 17085
rect 14553 17119 14611 17125
rect 14553 17085 14565 17119
rect 14599 17085 14611 17119
rect 14553 17079 14611 17085
rect 6963 17020 9076 17048
rect 9125 17051 9183 17057
rect 6963 17017 6975 17020
rect 6917 17011 6975 17017
rect 9125 17017 9137 17051
rect 9171 17048 9183 17051
rect 14292 17048 14320 17079
rect 14642 17076 14648 17128
rect 14700 17076 14706 17128
rect 14829 17119 14887 17125
rect 14829 17085 14841 17119
rect 14875 17116 14887 17119
rect 15289 17119 15347 17125
rect 15289 17116 15301 17119
rect 14875 17088 15301 17116
rect 14875 17085 14887 17088
rect 14829 17079 14887 17085
rect 15289 17085 15301 17088
rect 15335 17085 15347 17119
rect 15289 17079 15347 17085
rect 14458 17048 14464 17060
rect 9171 17020 9996 17048
rect 14292 17020 14464 17048
rect 9171 17017 9183 17020
rect 9125 17011 9183 17017
rect 9968 16992 9996 17020
rect 14458 17008 14464 17020
rect 14516 17048 14522 17060
rect 14844 17048 14872 17079
rect 16114 17076 16120 17128
rect 16172 17116 16178 17128
rect 16577 17119 16635 17125
rect 16577 17116 16589 17119
rect 16172 17088 16589 17116
rect 16172 17076 16178 17088
rect 16577 17085 16589 17088
rect 16623 17085 16635 17119
rect 16577 17079 16635 17085
rect 16666 17076 16672 17128
rect 16724 17076 16730 17128
rect 16758 17076 16764 17128
rect 16816 17116 16822 17128
rect 17037 17119 17095 17125
rect 17037 17116 17049 17119
rect 16816 17088 17049 17116
rect 16816 17076 16822 17088
rect 17037 17085 17049 17088
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 17313 17119 17371 17125
rect 17313 17085 17325 17119
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 14516 17020 14872 17048
rect 14516 17008 14522 17020
rect 15194 17008 15200 17060
rect 15252 17008 15258 17060
rect 15657 17051 15715 17057
rect 15657 17017 15669 17051
rect 15703 17048 15715 17051
rect 16850 17048 16856 17060
rect 15703 17020 16856 17048
rect 15703 17017 15715 17020
rect 15657 17011 15715 17017
rect 16850 17008 16856 17020
rect 16908 17008 16914 17060
rect 16945 17051 17003 17057
rect 16945 17017 16957 17051
rect 16991 17048 17003 17051
rect 17126 17048 17132 17060
rect 16991 17020 17132 17048
rect 16991 17017 17003 17020
rect 16945 17011 17003 17017
rect 17126 17008 17132 17020
rect 17184 17008 17190 17060
rect 5224 16952 5948 16980
rect 5224 16940 5230 16952
rect 6086 16940 6092 16992
rect 6144 16940 6150 16992
rect 9026 16983 9084 16989
rect 9026 16949 9038 16983
rect 9072 16980 9084 16983
rect 9766 16980 9772 16992
rect 9072 16952 9772 16980
rect 9072 16949 9084 16952
rect 9026 16943 9084 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 9950 16940 9956 16992
rect 10008 16940 10014 16992
rect 14369 16983 14427 16989
rect 14369 16949 14381 16983
rect 14415 16980 14427 16983
rect 14642 16980 14648 16992
rect 14415 16952 14648 16980
rect 14415 16949 14427 16952
rect 14369 16943 14427 16949
rect 14642 16940 14648 16952
rect 14700 16940 14706 16992
rect 16206 16940 16212 16992
rect 16264 16980 16270 16992
rect 16758 16980 16764 16992
rect 16264 16952 16764 16980
rect 16264 16940 16270 16952
rect 16758 16940 16764 16952
rect 16816 16980 16822 16992
rect 17328 16980 17356 17079
rect 17586 17076 17592 17128
rect 17644 17076 17650 17128
rect 17972 17116 18000 17215
rect 18046 17144 18052 17196
rect 18104 17184 18110 17196
rect 18104 17156 18828 17184
rect 18104 17144 18110 17156
rect 18325 17119 18383 17125
rect 18325 17116 18337 17119
rect 17972 17088 18337 17116
rect 18325 17085 18337 17088
rect 18371 17116 18383 17119
rect 18414 17116 18420 17128
rect 18371 17088 18420 17116
rect 18371 17085 18383 17088
rect 18325 17079 18383 17085
rect 18414 17076 18420 17088
rect 18472 17076 18478 17128
rect 18509 17119 18567 17125
rect 18509 17085 18521 17119
rect 18555 17116 18567 17119
rect 18598 17116 18604 17128
rect 18555 17088 18604 17116
rect 18555 17085 18567 17088
rect 18509 17079 18567 17085
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 18690 17076 18696 17128
rect 18748 17076 18754 17128
rect 18800 17116 18828 17156
rect 18949 17119 19007 17125
rect 18949 17116 18961 17119
rect 18800 17088 18961 17116
rect 18949 17085 18961 17088
rect 18995 17085 19007 17119
rect 18949 17079 19007 17085
rect 19518 17076 19524 17128
rect 19576 17116 19582 17128
rect 20824 17125 20852 17292
rect 22094 17280 22100 17292
rect 22152 17280 22158 17332
rect 22186 17280 22192 17332
rect 22244 17320 22250 17332
rect 22373 17323 22431 17329
rect 22373 17320 22385 17323
rect 22244 17292 22385 17320
rect 22244 17280 22250 17292
rect 22373 17289 22385 17292
rect 22419 17289 22431 17323
rect 22373 17283 22431 17289
rect 20717 17119 20775 17125
rect 20717 17116 20729 17119
rect 19576 17088 20729 17116
rect 19576 17076 19582 17088
rect 20717 17085 20729 17088
rect 20763 17116 20775 17119
rect 20809 17119 20867 17125
rect 20809 17116 20821 17119
rect 20763 17088 20821 17116
rect 20763 17085 20775 17088
rect 20717 17079 20775 17085
rect 20809 17085 20821 17088
rect 20855 17085 20867 17119
rect 21634 17116 21640 17128
rect 20809 17079 20867 17085
rect 21008 17088 21640 17116
rect 17402 17008 17408 17060
rect 17460 17048 17466 17060
rect 18708 17048 18736 17076
rect 17460 17020 18736 17048
rect 17460 17008 17466 17020
rect 19978 17008 19984 17060
rect 20036 17048 20042 17060
rect 20533 17051 20591 17057
rect 20533 17048 20545 17051
rect 20036 17020 20545 17048
rect 20036 17008 20042 17020
rect 20533 17017 20545 17020
rect 20579 17048 20591 17051
rect 21008 17048 21036 17088
rect 21634 17076 21640 17088
rect 21692 17076 21698 17128
rect 22186 17076 22192 17128
rect 22244 17116 22250 17128
rect 22649 17119 22707 17125
rect 22649 17116 22661 17119
rect 22244 17088 22661 17116
rect 22244 17076 22250 17088
rect 22649 17085 22661 17088
rect 22695 17085 22707 17119
rect 22649 17079 22707 17085
rect 20579 17020 21036 17048
rect 21076 17051 21134 17057
rect 20579 17017 20591 17020
rect 20533 17011 20591 17017
rect 21076 17017 21088 17051
rect 21122 17048 21134 17051
rect 21266 17048 21272 17060
rect 21122 17020 21272 17048
rect 21122 17017 21134 17020
rect 21076 17011 21134 17017
rect 21266 17008 21272 17020
rect 21324 17008 21330 17060
rect 16816 16952 17356 16980
rect 16816 16940 16822 16952
rect 17494 16940 17500 16992
rect 17552 16980 17558 16992
rect 19334 16980 19340 16992
rect 17552 16952 19340 16980
rect 17552 16940 17558 16952
rect 19334 16940 19340 16952
rect 19392 16940 19398 16992
rect 20070 16940 20076 16992
rect 20128 16940 20134 16992
rect 21726 16940 21732 16992
rect 21784 16980 21790 16992
rect 22189 16983 22247 16989
rect 22189 16980 22201 16983
rect 21784 16952 22201 16980
rect 21784 16940 21790 16952
rect 22189 16949 22201 16952
rect 22235 16949 22247 16983
rect 22189 16943 22247 16949
rect 552 16890 23368 16912
rect 552 16838 4322 16890
rect 4374 16838 4386 16890
rect 4438 16838 4450 16890
rect 4502 16838 4514 16890
rect 4566 16838 4578 16890
rect 4630 16838 23368 16890
rect 552 16816 23368 16838
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 5077 16779 5135 16785
rect 5077 16776 5089 16779
rect 4948 16748 5089 16776
rect 4948 16736 4954 16748
rect 5077 16745 5089 16748
rect 5123 16745 5135 16779
rect 5077 16739 5135 16745
rect 9490 16736 9496 16788
rect 9548 16736 9554 16788
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10061 16779 10119 16785
rect 10061 16776 10073 16779
rect 10008 16748 10073 16776
rect 10008 16736 10014 16748
rect 10061 16745 10073 16748
rect 10107 16745 10119 16779
rect 10061 16739 10119 16745
rect 14458 16736 14464 16788
rect 14516 16736 14522 16788
rect 16666 16736 16672 16788
rect 16724 16736 16730 16788
rect 18230 16736 18236 16788
rect 18288 16776 18294 16788
rect 19061 16779 19119 16785
rect 19061 16776 19073 16779
rect 18288 16748 19073 16776
rect 18288 16736 18294 16748
rect 19061 16745 19073 16748
rect 19107 16745 19119 16779
rect 19061 16739 19119 16745
rect 19334 16736 19340 16788
rect 19392 16776 19398 16788
rect 19392 16748 21220 16776
rect 19392 16736 19398 16748
rect 5442 16668 5448 16720
rect 5500 16708 5506 16720
rect 7466 16708 7472 16720
rect 5500 16680 6776 16708
rect 5500 16668 5506 16680
rect 4706 16600 4712 16652
rect 4764 16600 4770 16652
rect 4798 16600 4804 16652
rect 4856 16640 4862 16652
rect 4893 16643 4951 16649
rect 4893 16640 4905 16643
rect 4856 16612 4905 16640
rect 4856 16600 4862 16612
rect 4893 16609 4905 16612
rect 4939 16609 4951 16643
rect 4893 16603 4951 16609
rect 5902 16600 5908 16652
rect 5960 16640 5966 16652
rect 5997 16643 6055 16649
rect 5997 16640 6009 16643
rect 5960 16612 6009 16640
rect 5960 16600 5966 16612
rect 5997 16609 6009 16612
rect 6043 16609 6055 16643
rect 5997 16603 6055 16609
rect 4724 16572 4752 16600
rect 5534 16572 5540 16584
rect 4724 16544 5540 16572
rect 5534 16532 5540 16544
rect 5592 16572 5598 16584
rect 5810 16572 5816 16584
rect 5592 16544 5816 16572
rect 5592 16532 5598 16544
rect 5810 16532 5816 16544
rect 5868 16532 5874 16584
rect 6086 16532 6092 16584
rect 6144 16532 6150 16584
rect 6748 16581 6776 16680
rect 6840 16680 7472 16708
rect 6840 16649 6868 16680
rect 7466 16668 7472 16680
rect 7524 16668 7530 16720
rect 8570 16668 8576 16720
rect 8628 16708 8634 16720
rect 8628 16680 9628 16708
rect 8628 16668 8634 16680
rect 6825 16643 6883 16649
rect 6825 16609 6837 16643
rect 6871 16609 6883 16643
rect 6825 16603 6883 16609
rect 7098 16600 7104 16652
rect 7156 16600 7162 16652
rect 9306 16600 9312 16652
rect 9364 16600 9370 16652
rect 9600 16649 9628 16680
rect 9858 16668 9864 16720
rect 9916 16668 9922 16720
rect 15470 16708 15476 16720
rect 14936 16680 15476 16708
rect 9585 16643 9643 16649
rect 9585 16609 9597 16643
rect 9631 16609 9643 16643
rect 9585 16603 9643 16609
rect 9674 16600 9680 16652
rect 9732 16640 9738 16652
rect 9769 16643 9827 16649
rect 9769 16640 9781 16643
rect 9732 16612 9781 16640
rect 9732 16600 9738 16612
rect 9769 16609 9781 16612
rect 9815 16609 9827 16643
rect 9769 16603 9827 16609
rect 14645 16643 14703 16649
rect 14645 16609 14657 16643
rect 14691 16609 14703 16643
rect 14645 16603 14703 16609
rect 6733 16575 6791 16581
rect 6733 16541 6745 16575
rect 6779 16541 6791 16575
rect 14660 16572 14688 16603
rect 14826 16600 14832 16652
rect 14884 16600 14890 16652
rect 14936 16649 14964 16680
rect 15470 16668 15476 16680
rect 15528 16668 15534 16720
rect 15933 16711 15991 16717
rect 15933 16677 15945 16711
rect 15979 16708 15991 16711
rect 16206 16708 16212 16720
rect 15979 16680 16212 16708
rect 15979 16677 15991 16680
rect 15933 16671 15991 16677
rect 16206 16668 16212 16680
rect 16264 16708 16270 16720
rect 16684 16708 16712 16736
rect 16264 16680 17080 16708
rect 16264 16668 16270 16680
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16609 14979 16643
rect 14921 16603 14979 16609
rect 15010 16600 15016 16652
rect 15068 16600 15074 16652
rect 15197 16643 15255 16649
rect 15197 16609 15209 16643
rect 15243 16609 15255 16643
rect 15197 16603 15255 16609
rect 15105 16575 15163 16581
rect 15105 16572 15117 16575
rect 14660 16544 15117 16572
rect 6733 16535 6791 16541
rect 15105 16541 15117 16544
rect 15151 16541 15163 16575
rect 15105 16535 15163 16541
rect 6454 16464 6460 16516
rect 6512 16504 6518 16516
rect 7377 16507 7435 16513
rect 7377 16504 7389 16507
rect 6512 16476 7389 16504
rect 6512 16464 6518 16476
rect 7377 16473 7389 16476
rect 7423 16473 7435 16507
rect 7377 16467 7435 16473
rect 14458 16464 14464 16516
rect 14516 16504 14522 16516
rect 14918 16504 14924 16516
rect 14516 16476 14924 16504
rect 14516 16464 14522 16476
rect 14918 16464 14924 16476
rect 14976 16504 14982 16516
rect 15212 16504 15240 16603
rect 15378 16600 15384 16652
rect 15436 16640 15442 16652
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 15436 16612 15669 16640
rect 15436 16600 15442 16612
rect 15657 16609 15669 16612
rect 15703 16640 15715 16643
rect 15703 16612 16068 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16572 15807 16575
rect 15838 16572 15844 16584
rect 15795 16544 15844 16572
rect 15795 16541 15807 16544
rect 15749 16535 15807 16541
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 15930 16532 15936 16584
rect 15988 16532 15994 16584
rect 16040 16572 16068 16612
rect 16114 16600 16120 16652
rect 16172 16640 16178 16652
rect 16301 16643 16359 16649
rect 16301 16640 16313 16643
rect 16172 16612 16313 16640
rect 16172 16600 16178 16612
rect 16301 16609 16313 16612
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16640 16635 16643
rect 16666 16640 16672 16652
rect 16623 16612 16672 16640
rect 16623 16609 16635 16612
rect 16577 16603 16635 16609
rect 16666 16600 16672 16612
rect 16724 16600 16730 16652
rect 16758 16600 16764 16652
rect 16816 16640 16822 16652
rect 17052 16649 17080 16680
rect 17310 16668 17316 16720
rect 17368 16708 17374 16720
rect 20070 16708 20076 16720
rect 17368 16680 18736 16708
rect 17368 16668 17374 16680
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 16816 16612 16957 16640
rect 16816 16600 16822 16612
rect 16945 16609 16957 16612
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 17037 16643 17095 16649
rect 17037 16609 17049 16643
rect 17083 16609 17095 16643
rect 17037 16603 17095 16609
rect 17126 16600 17132 16652
rect 17184 16600 17190 16652
rect 18414 16600 18420 16652
rect 18472 16600 18478 16652
rect 18598 16600 18604 16652
rect 18656 16600 18662 16652
rect 18708 16640 18736 16680
rect 19076 16680 20076 16708
rect 19076 16649 19104 16680
rect 20070 16668 20076 16680
rect 20128 16668 20134 16720
rect 21192 16708 21220 16748
rect 21266 16736 21272 16788
rect 21324 16736 21330 16788
rect 22738 16708 22744 16720
rect 21192 16680 21404 16708
rect 19061 16643 19119 16649
rect 18708 16612 19012 16640
rect 16393 16575 16451 16581
rect 16393 16572 16405 16575
rect 16040 16544 16405 16572
rect 16393 16541 16405 16544
rect 16439 16541 16451 16575
rect 16393 16535 16451 16541
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 17310 16572 17316 16584
rect 16899 16544 17316 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 14976 16476 15240 16504
rect 15856 16504 15884 16532
rect 16485 16507 16543 16513
rect 16485 16504 16497 16507
rect 15856 16476 16497 16504
rect 14976 16464 14982 16476
rect 16485 16473 16497 16476
rect 16531 16473 16543 16507
rect 16485 16467 16543 16473
rect 16574 16464 16580 16516
rect 16632 16504 16638 16516
rect 16868 16504 16896 16535
rect 17310 16532 17316 16544
rect 17368 16532 17374 16584
rect 18984 16572 19012 16612
rect 19061 16609 19073 16643
rect 19107 16609 19119 16643
rect 19245 16643 19303 16649
rect 19245 16640 19257 16643
rect 19061 16603 19119 16609
rect 19168 16612 19257 16640
rect 19168 16572 19196 16612
rect 19245 16609 19257 16612
rect 19291 16640 19303 16643
rect 20530 16640 20536 16652
rect 19291 16612 20536 16640
rect 19291 16609 19303 16612
rect 19245 16603 19303 16609
rect 20530 16600 20536 16612
rect 20588 16600 20594 16652
rect 18984 16544 19196 16572
rect 21376 16572 21404 16680
rect 21468 16680 22744 16708
rect 21468 16649 21496 16680
rect 22738 16668 22744 16680
rect 22796 16668 22802 16720
rect 21453 16643 21511 16649
rect 21453 16609 21465 16643
rect 21499 16609 21511 16643
rect 21637 16643 21695 16649
rect 21637 16640 21649 16643
rect 21453 16603 21511 16609
rect 21560 16612 21649 16640
rect 21560 16572 21588 16612
rect 21637 16609 21649 16612
rect 21683 16609 21695 16643
rect 21637 16603 21695 16609
rect 21726 16600 21732 16652
rect 21784 16600 21790 16652
rect 21376 16544 21588 16572
rect 16632 16476 16896 16504
rect 16632 16464 16638 16476
rect 18322 16464 18328 16516
rect 18380 16504 18386 16516
rect 18417 16507 18475 16513
rect 18417 16504 18429 16507
rect 18380 16476 18429 16504
rect 18380 16464 18386 16476
rect 18417 16473 18429 16476
rect 18463 16473 18475 16507
rect 18417 16467 18475 16473
rect 6365 16439 6423 16445
rect 6365 16405 6377 16439
rect 6411 16436 6423 16439
rect 7190 16436 7196 16448
rect 6411 16408 7196 16436
rect 6411 16405 6423 16408
rect 6365 16399 6423 16405
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 7561 16439 7619 16445
rect 7561 16405 7573 16439
rect 7607 16436 7619 16439
rect 7742 16436 7748 16448
rect 7607 16408 7748 16436
rect 7607 16405 7619 16408
rect 7561 16399 7619 16405
rect 7742 16396 7748 16408
rect 7800 16396 7806 16448
rect 10042 16396 10048 16448
rect 10100 16396 10106 16448
rect 10226 16396 10232 16448
rect 10284 16396 10290 16448
rect 16114 16396 16120 16448
rect 16172 16396 16178 16448
rect 17034 16396 17040 16448
rect 17092 16436 17098 16448
rect 17313 16439 17371 16445
rect 17313 16436 17325 16439
rect 17092 16408 17325 16436
rect 17092 16396 17098 16408
rect 17313 16405 17325 16408
rect 17359 16405 17371 16439
rect 17313 16399 17371 16405
rect 552 16346 23368 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 23368 16346
rect 552 16272 23368 16294
rect 7098 16232 7104 16244
rect 6564 16204 7104 16232
rect 5074 16124 5080 16176
rect 5132 16164 5138 16176
rect 5169 16167 5227 16173
rect 5169 16164 5181 16167
rect 5132 16136 5181 16164
rect 5132 16124 5138 16136
rect 5169 16133 5181 16136
rect 5215 16133 5227 16167
rect 5169 16127 5227 16133
rect 6564 16105 6592 16204
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 7561 16235 7619 16241
rect 7561 16201 7573 16235
rect 7607 16232 7619 16235
rect 7607 16204 10732 16232
rect 7607 16201 7619 16204
rect 7561 16195 7619 16201
rect 6825 16167 6883 16173
rect 6825 16133 6837 16167
rect 6871 16164 6883 16167
rect 7466 16164 7472 16176
rect 6871 16136 7472 16164
rect 6871 16133 6883 16136
rect 6825 16127 6883 16133
rect 7466 16124 7472 16136
rect 7524 16164 7530 16176
rect 8941 16167 8999 16173
rect 7524 16136 8524 16164
rect 7524 16124 7530 16136
rect 6549 16099 6607 16105
rect 6549 16065 6561 16099
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 6914 16056 6920 16108
rect 6972 16056 6978 16108
rect 7190 16056 7196 16108
rect 7248 16096 7254 16108
rect 8496 16105 8524 16136
rect 8941 16133 8953 16167
rect 8987 16164 8999 16167
rect 8987 16136 9536 16164
rect 8987 16133 8999 16136
rect 8941 16127 8999 16133
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 7248 16068 7389 16096
rect 7248 16056 7254 16068
rect 7377 16065 7389 16068
rect 7423 16096 7435 16099
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7423 16068 7757 16096
rect 7423 16065 7435 16068
rect 7377 16059 7435 16065
rect 7745 16065 7757 16068
rect 7791 16065 7803 16099
rect 7745 16059 7803 16065
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 9030 16056 9036 16108
rect 9088 16096 9094 16108
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 9088 16068 9413 16096
rect 9088 16056 9094 16068
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 4893 16031 4951 16037
rect 4893 15997 4905 16031
rect 4939 16028 4951 16031
rect 5534 16028 5540 16040
rect 4939 16000 5540 16028
rect 4939 15997 4951 16000
rect 4893 15991 4951 15997
rect 5534 15988 5540 16000
rect 5592 16028 5598 16040
rect 6178 16028 6184 16040
rect 5592 16000 6184 16028
rect 5592 15988 5598 16000
rect 6178 15988 6184 16000
rect 6236 15988 6242 16040
rect 6454 15988 6460 16040
rect 6512 15988 6518 16040
rect 7285 16031 7343 16037
rect 7285 15997 7297 16031
rect 7331 16028 7343 16031
rect 7558 16028 7564 16040
rect 7331 16000 7564 16028
rect 7331 15997 7343 16000
rect 7285 15991 7343 15997
rect 7558 15988 7564 16000
rect 7616 15988 7622 16040
rect 7837 16031 7895 16037
rect 7837 15997 7849 16031
rect 7883 16028 7895 16031
rect 8570 16028 8576 16040
rect 7883 16000 8576 16028
rect 7883 15997 7895 16000
rect 7837 15991 7895 15997
rect 8570 15988 8576 16000
rect 8628 15988 8634 16040
rect 9508 16037 9536 16136
rect 10704 16096 10732 16204
rect 11808 16204 13216 16232
rect 11808 16105 11836 16204
rect 12986 16164 12992 16176
rect 11900 16136 12992 16164
rect 11793 16099 11851 16105
rect 11793 16096 11805 16099
rect 10704 16068 11805 16096
rect 11793 16065 11805 16068
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 9493 16031 9551 16037
rect 9493 15997 9505 16031
rect 9539 16028 9551 16031
rect 9674 16028 9680 16040
rect 9539 16000 9680 16028
rect 9539 15997 9551 16000
rect 9493 15991 9551 15997
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 10778 15988 10784 16040
rect 10836 15988 10842 16040
rect 11900 16037 11928 16136
rect 12986 16124 12992 16136
rect 13044 16124 13050 16176
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16096 12311 16099
rect 12621 16099 12679 16105
rect 12621 16096 12633 16099
rect 12299 16068 12633 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 12621 16065 12633 16068
rect 12667 16096 12679 16099
rect 12667 16068 13124 16096
rect 12667 16065 12679 16068
rect 12621 16059 12679 16065
rect 10874 16031 10932 16037
rect 10874 15997 10886 16031
rect 10920 15997 10932 16031
rect 10874 15991 10932 15997
rect 11885 16031 11943 16037
rect 11885 15997 11897 16031
rect 11931 15997 11943 16031
rect 11885 15991 11943 15997
rect 4798 15920 4804 15972
rect 4856 15960 4862 15972
rect 4985 15963 5043 15969
rect 4985 15960 4997 15963
rect 4856 15932 4997 15960
rect 4856 15920 4862 15932
rect 4985 15929 4997 15932
rect 5031 15929 5043 15963
rect 4985 15923 5043 15929
rect 5169 15963 5227 15969
rect 5169 15929 5181 15963
rect 5215 15960 5227 15963
rect 5626 15960 5632 15972
rect 5215 15932 5632 15960
rect 5215 15929 5227 15932
rect 5169 15923 5227 15929
rect 5626 15920 5632 15932
rect 5684 15920 5690 15972
rect 10318 15960 10324 15972
rect 9876 15932 10324 15960
rect 8110 15852 8116 15904
rect 8168 15892 8174 15904
rect 9876 15901 9904 15932
rect 10318 15920 10324 15932
rect 10376 15960 10382 15972
rect 10889 15960 10917 15991
rect 12526 15988 12532 16040
rect 12584 15988 12590 16040
rect 12986 15988 12992 16040
rect 13044 15988 13050 16040
rect 10376 15932 10917 15960
rect 10376 15920 10382 15932
rect 12250 15920 12256 15972
rect 12308 15960 12314 15972
rect 12544 15960 12572 15988
rect 13096 15960 13124 16068
rect 13188 16037 13216 16204
rect 14826 16192 14832 16244
rect 14884 16232 14890 16244
rect 15010 16232 15016 16244
rect 14884 16204 15016 16232
rect 14884 16192 14890 16204
rect 15010 16192 15016 16204
rect 15068 16232 15074 16244
rect 15289 16235 15347 16241
rect 15289 16232 15301 16235
rect 15068 16204 15301 16232
rect 15068 16192 15074 16204
rect 15289 16201 15301 16204
rect 15335 16201 15347 16235
rect 15289 16195 15347 16201
rect 15470 16192 15476 16244
rect 15528 16192 15534 16244
rect 16666 16192 16672 16244
rect 16724 16232 16730 16244
rect 16850 16232 16856 16244
rect 16724 16204 16856 16232
rect 16724 16192 16730 16204
rect 16850 16192 16856 16204
rect 16908 16232 16914 16244
rect 17221 16235 17279 16241
rect 17221 16232 17233 16235
rect 16908 16204 17233 16232
rect 16908 16192 16914 16204
rect 17221 16201 17233 16204
rect 17267 16232 17279 16235
rect 17494 16232 17500 16244
rect 17267 16204 17500 16232
rect 17267 16201 17279 16204
rect 17221 16195 17279 16201
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 19426 16192 19432 16244
rect 19484 16192 19490 16244
rect 20346 16192 20352 16244
rect 20404 16232 20410 16244
rect 21361 16235 21419 16241
rect 21361 16232 21373 16235
rect 20404 16204 21373 16232
rect 20404 16192 20410 16204
rect 13817 16167 13875 16173
rect 13817 16133 13829 16167
rect 13863 16164 13875 16167
rect 19981 16167 20039 16173
rect 19981 16164 19993 16167
rect 13863 16136 14964 16164
rect 13863 16133 13875 16136
rect 13817 16127 13875 16133
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16096 14611 16099
rect 14826 16096 14832 16108
rect 14599 16068 14832 16096
rect 14599 16065 14611 16068
rect 14553 16059 14611 16065
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 13173 16031 13231 16037
rect 13173 15997 13185 16031
rect 13219 15997 13231 16031
rect 13541 16031 13599 16037
rect 13541 16028 13553 16031
rect 13173 15991 13231 15997
rect 13280 16000 13553 16028
rect 13280 15960 13308 16000
rect 13541 15997 13553 16000
rect 13587 15997 13599 16031
rect 13541 15991 13599 15997
rect 14458 15988 14464 16040
rect 14516 16028 14522 16040
rect 14645 16031 14703 16037
rect 14645 16028 14657 16031
rect 14516 16000 14657 16028
rect 14516 15988 14522 16000
rect 14645 15997 14657 16000
rect 14691 15997 14703 16031
rect 14645 15991 14703 15997
rect 12308 15932 13032 15960
rect 13096 15932 13308 15960
rect 13357 15963 13415 15969
rect 12308 15920 12314 15932
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 8168 15864 8217 15892
rect 8168 15852 8174 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 8205 15855 8263 15861
rect 9861 15895 9919 15901
rect 9861 15861 9873 15895
rect 9907 15861 9919 15895
rect 9861 15855 9919 15861
rect 11149 15895 11207 15901
rect 11149 15861 11161 15895
rect 11195 15892 11207 15895
rect 11974 15892 11980 15904
rect 11195 15864 11980 15892
rect 11195 15861 11207 15864
rect 11149 15855 11207 15861
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 12894 15852 12900 15904
rect 12952 15852 12958 15904
rect 13004 15892 13032 15932
rect 13357 15929 13369 15963
rect 13403 15960 13415 15963
rect 13817 15963 13875 15969
rect 13817 15960 13829 15963
rect 13403 15932 13829 15960
rect 13403 15929 13415 15932
rect 13357 15923 13415 15929
rect 13817 15929 13829 15932
rect 13863 15929 13875 15963
rect 14660 15960 14688 15991
rect 14734 15988 14740 16040
rect 14792 16028 14798 16040
rect 14936 16037 14964 16136
rect 19352 16136 19993 16164
rect 15102 16056 15108 16108
rect 15160 16096 15166 16108
rect 15160 16068 15608 16096
rect 15160 16056 15166 16068
rect 15580 16037 15608 16068
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 14792 16000 14933 16028
rect 14792 15988 14798 16000
rect 14921 15997 14933 16000
rect 14967 15997 14979 16031
rect 15381 16031 15439 16037
rect 15381 16028 15393 16031
rect 14921 15991 14979 15997
rect 15028 16000 15393 16028
rect 15028 15960 15056 16000
rect 15381 15997 15393 16000
rect 15427 15997 15439 16031
rect 15381 15991 15439 15997
rect 15565 16031 15623 16037
rect 15565 15997 15577 16031
rect 15611 15997 15623 16031
rect 15565 15991 15623 15997
rect 16114 15988 16120 16040
rect 16172 15988 16178 16040
rect 16206 15988 16212 16040
rect 16264 16028 16270 16040
rect 16301 16031 16359 16037
rect 16301 16028 16313 16031
rect 16264 16000 16313 16028
rect 16264 15988 16270 16000
rect 16301 15997 16313 16000
rect 16347 15997 16359 16031
rect 16301 15991 16359 15997
rect 16482 15988 16488 16040
rect 16540 15988 16546 16040
rect 16942 15988 16948 16040
rect 17000 15988 17006 16040
rect 17034 15988 17040 16040
rect 17092 15988 17098 16040
rect 17313 16031 17371 16037
rect 17313 15997 17325 16031
rect 17359 16028 17371 16031
rect 17678 16028 17684 16040
rect 17359 16000 17684 16028
rect 17359 15997 17371 16000
rect 17313 15991 17371 15997
rect 17678 15988 17684 16000
rect 17736 15988 17742 16040
rect 18874 15988 18880 16040
rect 18932 16028 18938 16040
rect 19352 16037 19380 16136
rect 19981 16133 19993 16136
rect 20027 16133 20039 16167
rect 19981 16127 20039 16133
rect 19426 16056 19432 16108
rect 19484 16096 19490 16108
rect 19797 16099 19855 16105
rect 19797 16096 19809 16099
rect 19484 16068 19809 16096
rect 19484 16056 19490 16068
rect 19797 16065 19809 16068
rect 19843 16065 19855 16099
rect 19797 16059 19855 16065
rect 19904 16068 20116 16096
rect 19337 16031 19395 16037
rect 19337 16028 19349 16031
rect 18932 16000 19349 16028
rect 18932 15988 18938 16000
rect 19337 15997 19349 16000
rect 19383 15997 19395 16031
rect 19337 15991 19395 15997
rect 19518 15988 19524 16040
rect 19576 16028 19582 16040
rect 19904 16028 19932 16068
rect 20088 16040 20116 16068
rect 20548 16068 20944 16096
rect 19576 16000 19932 16028
rect 19576 15988 19582 16000
rect 20070 15988 20076 16040
rect 20128 15988 20134 16040
rect 20548 16037 20576 16068
rect 20916 16040 20944 16068
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 20809 16031 20867 16037
rect 20809 15997 20821 16031
rect 20855 15997 20867 16031
rect 20809 15991 20867 15997
rect 14660 15932 15056 15960
rect 15105 15963 15163 15969
rect 13817 15923 13875 15929
rect 15105 15929 15117 15963
rect 15151 15960 15163 15963
rect 15286 15960 15292 15972
rect 15151 15932 15292 15960
rect 15151 15929 15163 15932
rect 15105 15923 15163 15929
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 16393 15963 16451 15969
rect 16393 15929 16405 15963
rect 16439 15960 16451 15963
rect 17494 15960 17500 15972
rect 16439 15932 17500 15960
rect 16439 15929 16451 15932
rect 16393 15923 16451 15929
rect 17494 15920 17500 15932
rect 17552 15920 17558 15972
rect 20717 15963 20775 15969
rect 20717 15960 20729 15963
rect 19720 15932 20729 15960
rect 19720 15904 19748 15932
rect 20717 15929 20729 15932
rect 20763 15960 20775 15963
rect 20824 15960 20852 15991
rect 20898 15988 20904 16040
rect 20956 16028 20962 16040
rect 20993 16031 21051 16037
rect 20993 16028 21005 16031
rect 20956 16000 21005 16028
rect 20956 15988 20962 16000
rect 20993 15997 21005 16000
rect 21039 15997 21051 16031
rect 20993 15991 21051 15997
rect 20763 15932 20852 15960
rect 21192 15960 21220 16204
rect 21361 16201 21373 16204
rect 21407 16201 21419 16235
rect 21361 16195 21419 16201
rect 21821 16235 21879 16241
rect 21821 16201 21833 16235
rect 21867 16232 21879 16235
rect 22278 16232 22284 16244
rect 21867 16204 22284 16232
rect 21867 16201 21879 16204
rect 21821 16195 21879 16201
rect 21726 16164 21732 16176
rect 21284 16136 21732 16164
rect 21284 16037 21312 16136
rect 21726 16124 21732 16136
rect 21784 16124 21790 16176
rect 21545 16099 21603 16105
rect 21545 16065 21557 16099
rect 21591 16096 21603 16099
rect 21836 16096 21864 16195
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 21591 16068 21864 16096
rect 21591 16065 21603 16068
rect 21545 16059 21603 16065
rect 21269 16031 21327 16037
rect 21269 15997 21281 16031
rect 21315 15997 21327 16031
rect 21637 16031 21695 16037
rect 21637 16028 21649 16031
rect 21269 15991 21327 15997
rect 21468 16000 21649 16028
rect 21468 15972 21496 16000
rect 21637 15997 21649 16000
rect 21683 15997 21695 16031
rect 21637 15991 21695 15997
rect 21726 15988 21732 16040
rect 21784 15988 21790 16040
rect 22278 16028 22284 16040
rect 21836 16000 22284 16028
rect 21450 15960 21456 15972
rect 21192 15932 21456 15960
rect 20763 15929 20775 15932
rect 20717 15923 20775 15929
rect 21450 15920 21456 15932
rect 21508 15920 21514 15972
rect 21545 15963 21603 15969
rect 21545 15929 21557 15963
rect 21591 15960 21603 15963
rect 21836 15960 21864 16000
rect 22278 15988 22284 16000
rect 22336 15988 22342 16040
rect 22373 16031 22431 16037
rect 22373 15997 22385 16031
rect 22419 16028 22431 16031
rect 22646 16028 22652 16040
rect 22419 16000 22652 16028
rect 22419 15997 22431 16000
rect 22373 15991 22431 15997
rect 22646 15988 22652 16000
rect 22704 15988 22710 16040
rect 22094 15960 22100 15972
rect 21591 15932 21864 15960
rect 22020 15932 22100 15960
rect 21591 15929 21603 15932
rect 21545 15923 21603 15929
rect 13633 15895 13691 15901
rect 13633 15892 13645 15895
rect 13004 15864 13645 15892
rect 13633 15861 13645 15864
rect 13679 15861 13691 15895
rect 13633 15855 13691 15861
rect 14277 15895 14335 15901
rect 14277 15861 14289 15895
rect 14323 15892 14335 15895
rect 14366 15892 14372 15904
rect 14323 15864 14372 15892
rect 14323 15861 14335 15864
rect 14277 15855 14335 15861
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 16666 15852 16672 15904
rect 16724 15852 16730 15904
rect 16758 15852 16764 15904
rect 16816 15852 16822 15904
rect 19702 15852 19708 15904
rect 19760 15852 19766 15904
rect 19797 15895 19855 15901
rect 19797 15861 19809 15895
rect 19843 15892 19855 15895
rect 19886 15892 19892 15904
rect 19843 15864 19892 15892
rect 19843 15861 19855 15864
rect 19797 15855 19855 15861
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 20346 15852 20352 15904
rect 20404 15852 20410 15904
rect 20438 15852 20444 15904
rect 20496 15892 20502 15904
rect 22020 15901 22048 15932
rect 22094 15920 22100 15932
rect 22152 15960 22158 15972
rect 22189 15963 22247 15969
rect 22189 15960 22201 15963
rect 22152 15932 22201 15960
rect 22152 15920 22158 15932
rect 22189 15929 22201 15932
rect 22235 15929 22247 15963
rect 22189 15923 22247 15929
rect 20901 15895 20959 15901
rect 20901 15892 20913 15895
rect 20496 15864 20913 15892
rect 20496 15852 20502 15864
rect 20901 15861 20913 15864
rect 20947 15861 20959 15895
rect 20901 15855 20959 15861
rect 22005 15895 22063 15901
rect 22005 15861 22017 15895
rect 22051 15861 22063 15895
rect 22005 15855 22063 15861
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 22830 15892 22836 15904
rect 22612 15864 22836 15892
rect 22612 15852 22618 15864
rect 22830 15852 22836 15864
rect 22888 15852 22894 15904
rect 552 15802 23368 15824
rect 552 15750 4322 15802
rect 4374 15750 4386 15802
rect 4438 15750 4450 15802
rect 4502 15750 4514 15802
rect 4566 15750 4578 15802
rect 4630 15750 23368 15802
rect 552 15728 23368 15750
rect 5629 15691 5687 15697
rect 5629 15657 5641 15691
rect 5675 15657 5687 15691
rect 5629 15651 5687 15657
rect 4890 15580 4896 15632
rect 4948 15620 4954 15632
rect 5261 15623 5319 15629
rect 5261 15620 5273 15623
rect 4948 15592 5273 15620
rect 4948 15580 4954 15592
rect 5261 15589 5273 15592
rect 5307 15589 5319 15623
rect 5644 15620 5672 15651
rect 7558 15648 7564 15700
rect 7616 15648 7622 15700
rect 8481 15691 8539 15697
rect 8481 15657 8493 15691
rect 8527 15688 8539 15691
rect 10410 15688 10416 15700
rect 8527 15660 10416 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 10778 15688 10784 15700
rect 10520 15660 10784 15688
rect 6058 15623 6116 15629
rect 6058 15620 6070 15623
rect 5644 15592 6070 15620
rect 5261 15583 5319 15589
rect 6058 15589 6070 15592
rect 6104 15589 6116 15623
rect 6058 15583 6116 15589
rect 7742 15580 7748 15632
rect 7800 15580 7806 15632
rect 8036 15592 8616 15620
rect 5074 15512 5080 15564
rect 5132 15512 5138 15564
rect 5353 15555 5411 15561
rect 5353 15521 5365 15555
rect 5399 15521 5411 15555
rect 5353 15515 5411 15521
rect 5445 15555 5503 15561
rect 5445 15521 5457 15555
rect 5491 15552 5503 15555
rect 5626 15552 5632 15564
rect 5491 15524 5632 15552
rect 5491 15521 5503 15524
rect 5445 15515 5503 15521
rect 5368 15348 5396 15515
rect 5626 15512 5632 15524
rect 5684 15552 5690 15564
rect 6362 15552 6368 15564
rect 5684 15524 6368 15552
rect 5684 15512 5690 15524
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 7466 15512 7472 15564
rect 7524 15512 7530 15564
rect 5810 15444 5816 15496
rect 5868 15444 5874 15496
rect 8036 15493 8064 15592
rect 8110 15512 8116 15564
rect 8168 15512 8174 15564
rect 8588 15561 8616 15592
rect 8573 15555 8631 15561
rect 8573 15521 8585 15555
rect 8619 15521 8631 15555
rect 8573 15515 8631 15521
rect 8666 15555 8724 15561
rect 8666 15521 8678 15555
rect 8712 15521 8724 15555
rect 8666 15515 8724 15521
rect 8021 15487 8079 15493
rect 8021 15453 8033 15487
rect 8067 15453 8079 15487
rect 8128 15484 8156 15512
rect 8680 15484 8708 15515
rect 9030 15512 9036 15564
rect 9088 15552 9094 15564
rect 9585 15555 9643 15561
rect 9585 15552 9597 15555
rect 9088 15524 9597 15552
rect 9088 15512 9094 15524
rect 9585 15521 9597 15524
rect 9631 15521 9643 15555
rect 9585 15515 9643 15521
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 9732 15524 9777 15552
rect 9732 15512 9738 15524
rect 10318 15512 10324 15564
rect 10376 15512 10382 15564
rect 10520 15561 10548 15660
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 12250 15688 12256 15700
rect 11256 15660 12256 15688
rect 11256 15561 11284 15660
rect 12250 15648 12256 15660
rect 12308 15648 12314 15700
rect 12406 15660 12664 15688
rect 11330 15580 11336 15632
rect 11388 15620 11394 15632
rect 12406 15620 12434 15660
rect 11388 15592 12434 15620
rect 11388 15580 11394 15592
rect 10505 15555 10563 15561
rect 10505 15521 10517 15555
rect 10551 15521 10563 15555
rect 10505 15515 10563 15521
rect 11241 15555 11299 15561
rect 11241 15521 11253 15555
rect 11287 15521 11299 15555
rect 11241 15515 11299 15521
rect 11514 15512 11520 15564
rect 11572 15552 11578 15564
rect 11701 15555 11759 15561
rect 11701 15552 11713 15555
rect 11572 15524 11713 15552
rect 11572 15512 11578 15524
rect 11701 15521 11713 15524
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 11882 15512 11888 15564
rect 11940 15512 11946 15564
rect 11974 15512 11980 15564
rect 12032 15512 12038 15564
rect 12069 15555 12127 15561
rect 12069 15521 12081 15555
rect 12115 15521 12127 15555
rect 12069 15515 12127 15521
rect 8128 15456 8708 15484
rect 9953 15487 10011 15493
rect 8021 15447 8079 15453
rect 9953 15453 9965 15487
rect 9999 15484 10011 15487
rect 10336 15484 10364 15512
rect 10413 15487 10471 15493
rect 10413 15484 10425 15487
rect 9999 15456 10272 15484
rect 10336 15456 10425 15484
rect 9999 15453 10011 15456
rect 9953 15447 10011 15453
rect 7745 15419 7803 15425
rect 7745 15385 7757 15419
rect 7791 15416 7803 15419
rect 8036 15416 8064 15447
rect 7791 15388 8064 15416
rect 7791 15385 7803 15388
rect 7745 15379 7803 15385
rect 10134 15376 10140 15428
rect 10192 15376 10198 15428
rect 10244 15416 10272 15456
rect 10413 15453 10425 15456
rect 10459 15453 10471 15487
rect 10413 15447 10471 15453
rect 10686 15444 10692 15496
rect 10744 15484 10750 15496
rect 11149 15487 11207 15493
rect 11149 15484 11161 15487
rect 10744 15456 11161 15484
rect 10744 15444 10750 15456
rect 11149 15453 11161 15456
rect 11195 15484 11207 15487
rect 12084 15484 12112 15515
rect 12250 15512 12256 15564
rect 12308 15512 12314 15564
rect 12526 15552 12532 15564
rect 12406 15524 12532 15552
rect 11195 15456 12112 15484
rect 12161 15487 12219 15493
rect 11195 15453 11207 15456
rect 11149 15447 11207 15453
rect 12161 15453 12173 15487
rect 12207 15484 12219 15487
rect 12406 15484 12434 15524
rect 12526 15512 12532 15524
rect 12584 15512 12590 15564
rect 12636 15561 12664 15660
rect 17494 15648 17500 15700
rect 17552 15648 17558 15700
rect 20283 15691 20341 15697
rect 20283 15657 20295 15691
rect 20329 15688 20341 15691
rect 20438 15688 20444 15700
rect 20329 15660 20444 15688
rect 20329 15657 20341 15660
rect 20283 15651 20341 15657
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 15286 15620 15292 15632
rect 14568 15592 15292 15620
rect 12621 15555 12679 15561
rect 12621 15521 12633 15555
rect 12667 15552 12679 15555
rect 12710 15552 12716 15564
rect 12667 15524 12716 15552
rect 12667 15521 12679 15524
rect 12621 15515 12679 15521
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 12805 15555 12863 15561
rect 12805 15521 12817 15555
rect 12851 15552 12863 15555
rect 12894 15552 12900 15564
rect 12851 15524 12900 15552
rect 12851 15521 12863 15524
rect 12805 15515 12863 15521
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 14568 15561 14596 15592
rect 15286 15580 15292 15592
rect 15344 15580 15350 15632
rect 16384 15623 16442 15629
rect 16384 15589 16396 15623
rect 16430 15620 16442 15623
rect 16666 15620 16672 15632
rect 16430 15592 16672 15620
rect 16430 15589 16442 15592
rect 16384 15583 16442 15589
rect 16666 15580 16672 15592
rect 16724 15580 16730 15632
rect 20073 15623 20131 15629
rect 20073 15589 20085 15623
rect 20119 15620 20131 15623
rect 20898 15620 20904 15632
rect 20119 15592 20904 15620
rect 20119 15589 20131 15592
rect 20073 15583 20131 15589
rect 20898 15580 20904 15592
rect 20956 15580 20962 15632
rect 14553 15555 14611 15561
rect 14553 15521 14565 15555
rect 14599 15521 14611 15555
rect 14553 15515 14611 15521
rect 14734 15512 14740 15564
rect 14792 15512 14798 15564
rect 17402 15552 17408 15564
rect 16132 15524 17408 15552
rect 16132 15496 16160 15524
rect 17402 15512 17408 15524
rect 17460 15512 17466 15564
rect 17678 15512 17684 15564
rect 17736 15512 17742 15564
rect 17862 15512 17868 15564
rect 17920 15512 17926 15564
rect 18785 15555 18843 15561
rect 18785 15521 18797 15555
rect 18831 15552 18843 15555
rect 19518 15552 19524 15564
rect 18831 15524 19524 15552
rect 18831 15521 18843 15524
rect 18785 15515 18843 15521
rect 19518 15512 19524 15524
rect 19576 15512 19582 15564
rect 19702 15512 19708 15564
rect 19760 15512 19766 15564
rect 19886 15512 19892 15564
rect 19944 15512 19950 15564
rect 20530 15512 20536 15564
rect 20588 15512 20594 15564
rect 20809 15555 20867 15561
rect 20809 15552 20821 15555
rect 20732 15524 20821 15552
rect 12207 15456 12434 15484
rect 12207 15453 12219 15456
rect 12161 15447 12219 15453
rect 13814 15444 13820 15496
rect 13872 15444 13878 15496
rect 16114 15444 16120 15496
rect 16172 15444 16178 15496
rect 18874 15444 18880 15496
rect 18932 15444 18938 15496
rect 20622 15444 20628 15496
rect 20680 15444 20686 15496
rect 11882 15416 11888 15428
rect 10244 15388 11888 15416
rect 11882 15376 11888 15388
rect 11940 15376 11946 15428
rect 20441 15419 20499 15425
rect 20441 15385 20453 15419
rect 20487 15416 20499 15419
rect 20732 15416 20760 15524
rect 20809 15521 20821 15524
rect 20855 15521 20867 15555
rect 20809 15515 20867 15521
rect 21637 15555 21695 15561
rect 21637 15521 21649 15555
rect 21683 15552 21695 15555
rect 21726 15552 21732 15564
rect 21683 15524 21732 15552
rect 21683 15521 21695 15524
rect 21637 15515 21695 15521
rect 21726 15512 21732 15524
rect 21784 15512 21790 15564
rect 22281 15555 22339 15561
rect 22281 15521 22293 15555
rect 22327 15552 22339 15555
rect 22646 15552 22652 15564
rect 22327 15524 22652 15552
rect 22327 15521 22339 15524
rect 22281 15515 22339 15521
rect 22646 15512 22652 15524
rect 22704 15512 22710 15564
rect 21450 15444 21456 15496
rect 21508 15484 21514 15496
rect 21545 15487 21603 15493
rect 21545 15484 21557 15487
rect 21508 15456 21557 15484
rect 21508 15444 21514 15456
rect 21545 15453 21557 15456
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 22189 15487 22247 15493
rect 22189 15484 22201 15487
rect 22152 15456 22201 15484
rect 22152 15444 22158 15456
rect 22189 15453 22201 15456
rect 22235 15453 22247 15487
rect 22189 15447 22247 15453
rect 20487 15388 20760 15416
rect 20993 15419 21051 15425
rect 20487 15385 20499 15388
rect 20441 15379 20499 15385
rect 20993 15385 21005 15419
rect 21039 15416 21051 15419
rect 22002 15416 22008 15428
rect 21039 15388 22008 15416
rect 21039 15385 21051 15388
rect 20993 15379 21051 15385
rect 22002 15376 22008 15388
rect 22060 15376 22066 15428
rect 6546 15348 6552 15360
rect 5368 15320 6552 15348
rect 6546 15308 6552 15320
rect 6604 15348 6610 15360
rect 7193 15351 7251 15357
rect 7193 15348 7205 15351
rect 6604 15320 7205 15348
rect 6604 15308 6610 15320
rect 7193 15317 7205 15320
rect 7239 15317 7251 15351
rect 7193 15311 7251 15317
rect 8757 15351 8815 15357
rect 8757 15317 8769 15351
rect 8803 15348 8815 15351
rect 11330 15348 11336 15360
rect 8803 15320 11336 15348
rect 8803 15317 8815 15320
rect 8757 15311 8815 15317
rect 11330 15308 11336 15320
rect 11388 15308 11394 15360
rect 11514 15308 11520 15360
rect 11572 15308 11578 15360
rect 11606 15308 11612 15360
rect 11664 15348 11670 15360
rect 11701 15351 11759 15357
rect 11701 15348 11713 15351
rect 11664 15320 11713 15348
rect 11664 15308 11670 15320
rect 11701 15317 11713 15320
rect 11747 15317 11759 15351
rect 11701 15311 11759 15317
rect 12989 15351 13047 15357
rect 12989 15317 13001 15351
rect 13035 15348 13047 15351
rect 13538 15348 13544 15360
rect 13035 15320 13544 15348
rect 13035 15317 13047 15320
rect 12989 15311 13047 15317
rect 13538 15308 13544 15320
rect 13596 15308 13602 15360
rect 17770 15308 17776 15360
rect 17828 15308 17834 15360
rect 18414 15308 18420 15360
rect 18472 15308 18478 15360
rect 19794 15308 19800 15360
rect 19852 15308 19858 15360
rect 20257 15351 20315 15357
rect 20257 15317 20269 15351
rect 20303 15348 20315 15351
rect 20346 15348 20352 15360
rect 20303 15320 20352 15348
rect 20303 15317 20315 15320
rect 20257 15311 20315 15317
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 20622 15308 20628 15360
rect 20680 15308 20686 15360
rect 21266 15308 21272 15360
rect 21324 15308 21330 15360
rect 21913 15351 21971 15357
rect 21913 15317 21925 15351
rect 21959 15348 21971 15351
rect 22370 15348 22376 15360
rect 21959 15320 22376 15348
rect 21959 15317 21971 15320
rect 21913 15311 21971 15317
rect 22370 15308 22376 15320
rect 22428 15308 22434 15360
rect 552 15258 23368 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 23368 15258
rect 552 15184 23368 15206
rect 10962 15104 10968 15156
rect 11020 15104 11026 15156
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 12032 15116 12173 15144
rect 12032 15104 12038 15116
rect 12161 15113 12173 15116
rect 12207 15113 12219 15147
rect 12161 15107 12219 15113
rect 12526 15104 12532 15156
rect 12584 15144 12590 15156
rect 12897 15147 12955 15153
rect 12897 15144 12909 15147
rect 12584 15116 12909 15144
rect 12584 15104 12590 15116
rect 12897 15113 12909 15116
rect 12943 15113 12955 15147
rect 12897 15107 12955 15113
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 13909 15147 13967 15153
rect 13909 15144 13921 15147
rect 13872 15116 13921 15144
rect 13872 15104 13878 15116
rect 13909 15113 13921 15116
rect 13955 15113 13967 15147
rect 13909 15107 13967 15113
rect 9398 15076 9404 15088
rect 8956 15048 9404 15076
rect 8956 15017 8984 15048
rect 9398 15036 9404 15048
rect 9456 15036 9462 15088
rect 8941 15011 8999 15017
rect 8941 14977 8953 15011
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 9214 14968 9220 15020
rect 9272 14968 9278 15020
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 11992 15008 12020 15104
rect 13078 15036 13084 15088
rect 13136 15076 13142 15088
rect 13136 15048 13860 15076
rect 13136 15036 13142 15048
rect 13832 15017 13860 15048
rect 9824 14980 10456 15008
rect 9824 14968 9830 14980
rect 8849 14943 8907 14949
rect 8849 14909 8861 14943
rect 8895 14940 8907 14943
rect 9122 14940 9128 14952
rect 8895 14912 9128 14940
rect 8895 14909 8907 14912
rect 8849 14903 8907 14909
rect 9122 14900 9128 14912
rect 9180 14940 9186 14952
rect 9309 14943 9367 14949
rect 9309 14940 9321 14943
rect 9180 14912 9321 14940
rect 9180 14900 9186 14912
rect 9309 14909 9321 14912
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 9398 14900 9404 14952
rect 9456 14940 9462 14952
rect 9861 14943 9919 14949
rect 9456 14912 9501 14940
rect 9456 14900 9462 14912
rect 9861 14909 9873 14943
rect 9907 14940 9919 14943
rect 9950 14940 9956 14952
rect 9907 14912 9956 14940
rect 9907 14909 9919 14912
rect 9861 14903 9919 14909
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 10045 14943 10103 14949
rect 10045 14909 10057 14943
rect 10091 14940 10103 14943
rect 10318 14940 10324 14952
rect 10091 14912 10324 14940
rect 10091 14909 10103 14912
rect 10045 14903 10103 14909
rect 10318 14900 10324 14912
rect 10376 14900 10382 14952
rect 10428 14949 10456 14980
rect 11440 14980 12020 15008
rect 13817 15011 13875 15017
rect 11440 14949 11468 14980
rect 13817 14977 13829 15011
rect 13863 14977 13875 15011
rect 13924 15008 13952 15107
rect 14642 15104 14648 15156
rect 14700 15144 14706 15156
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 14700 15116 14933 15144
rect 14700 15104 14706 15116
rect 14921 15113 14933 15116
rect 14967 15113 14979 15147
rect 14921 15107 14979 15113
rect 17678 15104 17684 15156
rect 17736 15144 17742 15156
rect 17865 15147 17923 15153
rect 17865 15144 17877 15147
rect 17736 15116 17877 15144
rect 17736 15104 17742 15116
rect 17865 15113 17877 15116
rect 17911 15113 17923 15147
rect 17865 15107 17923 15113
rect 18325 15147 18383 15153
rect 18325 15113 18337 15147
rect 18371 15144 18383 15147
rect 18874 15144 18880 15156
rect 18371 15116 18880 15144
rect 18371 15113 18383 15116
rect 18325 15107 18383 15113
rect 14277 15079 14335 15085
rect 14277 15045 14289 15079
rect 14323 15076 14335 15079
rect 15194 15076 15200 15088
rect 14323 15048 15200 15076
rect 14323 15045 14335 15048
rect 14277 15039 14335 15045
rect 15194 15036 15200 15048
rect 15252 15036 15258 15088
rect 14090 15008 14096 15020
rect 13924 14980 14096 15008
rect 13817 14971 13875 14977
rect 14090 14968 14096 14980
rect 14148 15008 14154 15020
rect 14148 14980 14504 15008
rect 14148 14968 14154 14980
rect 10413 14943 10471 14949
rect 10413 14909 10425 14943
rect 10459 14909 10471 14943
rect 10413 14903 10471 14909
rect 11425 14943 11483 14949
rect 11425 14909 11437 14943
rect 11471 14909 11483 14943
rect 11425 14903 11483 14909
rect 11514 14900 11520 14952
rect 11572 14940 11578 14952
rect 11701 14943 11759 14949
rect 11701 14940 11713 14943
rect 11572 14912 11713 14940
rect 11572 14900 11578 14912
rect 11701 14909 11713 14912
rect 11747 14940 11759 14943
rect 11747 14912 12112 14940
rect 11747 14909 11759 14912
rect 11701 14903 11759 14909
rect 10134 14832 10140 14884
rect 10192 14872 10198 14884
rect 10229 14875 10287 14881
rect 10229 14872 10241 14875
rect 10192 14844 10241 14872
rect 10192 14832 10198 14844
rect 10229 14841 10241 14844
rect 10275 14841 10287 14875
rect 10781 14875 10839 14881
rect 10229 14835 10287 14841
rect 10520 14844 10732 14872
rect 9677 14807 9735 14813
rect 9677 14773 9689 14807
rect 9723 14804 9735 14807
rect 9766 14804 9772 14816
rect 9723 14776 9772 14804
rect 9723 14773 9735 14776
rect 9677 14767 9735 14773
rect 9766 14764 9772 14776
rect 9824 14764 9830 14816
rect 10045 14807 10103 14813
rect 10045 14773 10057 14807
rect 10091 14804 10103 14807
rect 10520 14804 10548 14844
rect 10091 14776 10548 14804
rect 10091 14773 10103 14776
rect 10045 14767 10103 14773
rect 10594 14764 10600 14816
rect 10652 14764 10658 14816
rect 10704 14804 10732 14844
rect 10781 14841 10793 14875
rect 10827 14872 10839 14875
rect 11330 14872 11336 14884
rect 10827 14844 11336 14872
rect 10827 14841 10839 14844
rect 10781 14835 10839 14841
rect 11330 14832 11336 14844
rect 11388 14832 11394 14884
rect 11977 14875 12035 14881
rect 11977 14872 11989 14875
rect 11808 14844 11989 14872
rect 11808 14816 11836 14844
rect 11977 14841 11989 14844
rect 12023 14841 12035 14875
rect 12084 14872 12112 14912
rect 13538 14900 13544 14952
rect 13596 14940 13602 14952
rect 14001 14943 14059 14949
rect 13596 14912 13952 14940
rect 13596 14900 13602 14912
rect 12177 14875 12235 14881
rect 12177 14872 12189 14875
rect 12084 14844 12189 14872
rect 11977 14835 12035 14841
rect 12177 14841 12189 14844
rect 12223 14841 12235 14875
rect 12177 14835 12235 14841
rect 12710 14832 12716 14884
rect 12768 14832 12774 14884
rect 12894 14832 12900 14884
rect 12952 14881 12958 14884
rect 12952 14875 12971 14881
rect 12959 14841 12971 14875
rect 13924 14872 13952 14912
rect 14001 14909 14013 14943
rect 14047 14940 14059 14943
rect 14366 14940 14372 14952
rect 14047 14912 14372 14940
rect 14047 14909 14059 14912
rect 14001 14903 14059 14909
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 14476 14949 14504 14980
rect 14461 14943 14519 14949
rect 14461 14909 14473 14943
rect 14507 14909 14519 14943
rect 14461 14903 14519 14909
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14909 14703 14943
rect 14645 14903 14703 14909
rect 14737 14943 14795 14949
rect 14737 14909 14749 14943
rect 14783 14909 14795 14943
rect 14737 14903 14795 14909
rect 14660 14872 14688 14903
rect 12952 14835 12971 14841
rect 13004 14844 13676 14872
rect 13924 14844 14688 14872
rect 12952 14832 12958 14835
rect 10870 14804 10876 14816
rect 10704 14776 10876 14804
rect 10870 14764 10876 14776
rect 10928 14804 10934 14816
rect 10981 14807 11039 14813
rect 10981 14804 10993 14807
rect 10928 14776 10993 14804
rect 10928 14764 10934 14776
rect 10981 14773 10993 14776
rect 11027 14773 11039 14807
rect 10981 14767 11039 14773
rect 11149 14807 11207 14813
rect 11149 14773 11161 14807
rect 11195 14804 11207 14807
rect 11422 14804 11428 14816
rect 11195 14776 11428 14804
rect 11195 14773 11207 14776
rect 11149 14767 11207 14773
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 11517 14807 11575 14813
rect 11517 14773 11529 14807
rect 11563 14804 11575 14807
rect 11790 14804 11796 14816
rect 11563 14776 11796 14804
rect 11563 14773 11575 14776
rect 11517 14767 11575 14773
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 11882 14764 11888 14816
rect 11940 14764 11946 14816
rect 12342 14764 12348 14816
rect 12400 14804 12406 14816
rect 13004 14804 13032 14844
rect 13648 14813 13676 14844
rect 12400 14776 13032 14804
rect 13633 14807 13691 14813
rect 12400 14764 12406 14776
rect 13633 14773 13645 14807
rect 13679 14773 13691 14807
rect 13633 14767 13691 14773
rect 14642 14764 14648 14816
rect 14700 14804 14706 14816
rect 14752 14804 14780 14903
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 16114 14940 16120 14952
rect 15528 14912 16120 14940
rect 15528 14900 15534 14912
rect 16114 14900 16120 14912
rect 16172 14940 16178 14952
rect 16758 14949 16764 14952
rect 16485 14943 16543 14949
rect 16485 14940 16497 14943
rect 16172 14912 16497 14940
rect 16172 14900 16178 14912
rect 16485 14909 16497 14912
rect 16531 14909 16543 14943
rect 16752 14940 16764 14949
rect 16719 14912 16764 14940
rect 16485 14903 16543 14909
rect 16752 14903 16764 14912
rect 16758 14900 16764 14903
rect 16816 14900 16822 14952
rect 17880 14940 17908 15107
rect 18141 14943 18199 14949
rect 18141 14940 18153 14943
rect 17880 14912 18153 14940
rect 18141 14909 18153 14912
rect 18187 14909 18199 14943
rect 18141 14903 18199 14909
rect 17862 14832 17868 14884
rect 17920 14872 17926 14884
rect 17957 14875 18015 14881
rect 17957 14872 17969 14875
rect 17920 14844 17969 14872
rect 17920 14832 17926 14844
rect 17957 14841 17969 14844
rect 18003 14841 18015 14875
rect 17957 14835 18015 14841
rect 14700 14776 14780 14804
rect 14700 14764 14706 14776
rect 17586 14764 17592 14816
rect 17644 14804 17650 14816
rect 18340 14804 18368 15107
rect 18874 15104 18880 15116
rect 18932 15144 18938 15156
rect 19242 15144 19248 15156
rect 18932 15116 19248 15144
rect 18932 15104 18938 15116
rect 19242 15104 19248 15116
rect 19300 15104 19306 15156
rect 20622 15104 20628 15156
rect 20680 15144 20686 15156
rect 20717 15147 20775 15153
rect 20717 15144 20729 15147
rect 20680 15116 20729 15144
rect 20680 15104 20686 15116
rect 20717 15113 20729 15116
rect 20763 15113 20775 15147
rect 20717 15107 20775 15113
rect 21821 15079 21879 15085
rect 21821 15045 21833 15079
rect 21867 15076 21879 15079
rect 22097 15079 22155 15085
rect 22097 15076 22109 15079
rect 21867 15048 22109 15076
rect 21867 15045 21879 15048
rect 21821 15039 21879 15045
rect 22097 15045 22109 15048
rect 22143 15045 22155 15079
rect 22097 15039 22155 15045
rect 19794 14968 19800 15020
rect 19852 14968 19858 15020
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 15008 20315 15011
rect 20714 15008 20720 15020
rect 20303 14980 20720 15008
rect 20303 14977 20315 14980
rect 20257 14971 20315 14977
rect 20714 14968 20720 14980
rect 20772 14968 20778 15020
rect 21266 14968 21272 15020
rect 21324 15008 21330 15020
rect 21361 15011 21419 15017
rect 21361 15008 21373 15011
rect 21324 14980 21373 15008
rect 21324 14968 21330 14980
rect 21361 14977 21373 14980
rect 21407 14977 21419 15011
rect 21361 14971 21419 14977
rect 21913 15011 21971 15017
rect 21913 14977 21925 15011
rect 21959 15008 21971 15011
rect 22465 15011 22523 15017
rect 22465 15008 22477 15011
rect 21959 14980 22477 15008
rect 21959 14977 21971 14980
rect 21913 14971 21971 14977
rect 22465 14977 22477 14980
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 19886 14900 19892 14952
rect 19944 14900 19950 14952
rect 20438 14900 20444 14952
rect 20496 14900 20502 14952
rect 21450 14900 21456 14952
rect 21508 14900 21514 14952
rect 22002 14900 22008 14952
rect 22060 14900 22066 14952
rect 22370 14900 22376 14952
rect 22428 14940 22434 14952
rect 22649 14943 22707 14949
rect 22649 14940 22661 14943
rect 22428 14912 22661 14940
rect 22428 14900 22434 14912
rect 22649 14909 22661 14912
rect 22695 14909 22707 14943
rect 22649 14903 22707 14909
rect 22741 14943 22799 14949
rect 22741 14909 22753 14943
rect 22787 14909 22799 14943
rect 22741 14903 22799 14909
rect 18690 14832 18696 14884
rect 18748 14832 18754 14884
rect 18874 14832 18880 14884
rect 18932 14832 18938 14884
rect 20346 14832 20352 14884
rect 20404 14872 20410 14884
rect 20533 14875 20591 14881
rect 20533 14872 20545 14875
rect 20404 14844 20545 14872
rect 20404 14832 20410 14844
rect 20533 14841 20545 14844
rect 20579 14841 20591 14875
rect 20533 14835 20591 14841
rect 20717 14875 20775 14881
rect 20717 14841 20729 14875
rect 20763 14872 20775 14875
rect 20898 14872 20904 14884
rect 20763 14844 20904 14872
rect 20763 14841 20775 14844
rect 20717 14835 20775 14841
rect 20898 14832 20904 14844
rect 20956 14832 20962 14884
rect 22281 14875 22339 14881
rect 22281 14841 22293 14875
rect 22327 14872 22339 14875
rect 22554 14872 22560 14884
rect 22327 14844 22560 14872
rect 22327 14841 22339 14844
rect 22281 14835 22339 14841
rect 22554 14832 22560 14844
rect 22612 14872 22618 14884
rect 22756 14872 22784 14903
rect 22612 14844 22784 14872
rect 22612 14832 22618 14844
rect 17644 14776 18368 14804
rect 17644 14764 17650 14776
rect 19058 14764 19064 14816
rect 19116 14764 19122 14816
rect 22462 14764 22468 14816
rect 22520 14764 22526 14816
rect 552 14714 23368 14736
rect 552 14662 4322 14714
rect 4374 14662 4386 14714
rect 4438 14662 4450 14714
rect 4502 14662 4514 14714
rect 4566 14662 4578 14714
rect 4630 14662 23368 14714
rect 552 14640 23368 14662
rect 6178 14560 6184 14612
rect 6236 14560 6242 14612
rect 10134 14600 10140 14612
rect 9692 14572 10140 14600
rect 9692 14544 9720 14572
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 10962 14600 10968 14612
rect 10643 14572 10968 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 10962 14560 10968 14572
rect 11020 14600 11026 14612
rect 11020 14572 11284 14600
rect 11020 14560 11026 14572
rect 9674 14492 9680 14544
rect 9732 14492 9738 14544
rect 11256 14541 11284 14572
rect 11882 14560 11888 14612
rect 11940 14600 11946 14612
rect 12897 14603 12955 14609
rect 12897 14600 12909 14603
rect 11940 14572 12909 14600
rect 11940 14560 11946 14572
rect 12897 14569 12909 14572
rect 12943 14600 12955 14603
rect 13170 14600 13176 14612
rect 12943 14572 13176 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 14366 14560 14372 14612
rect 14424 14600 14430 14612
rect 14527 14603 14585 14609
rect 14527 14600 14539 14603
rect 14424 14572 14539 14600
rect 14424 14560 14430 14572
rect 14527 14569 14539 14572
rect 14573 14600 14585 14603
rect 14573 14572 14872 14600
rect 14573 14569 14585 14572
rect 14527 14563 14585 14569
rect 9861 14535 9919 14541
rect 9861 14501 9873 14535
rect 9907 14532 9919 14535
rect 11241 14535 11299 14541
rect 9907 14504 10272 14532
rect 9907 14501 9919 14504
rect 9861 14495 9919 14501
rect 10244 14476 10272 14504
rect 11241 14501 11253 14535
rect 11287 14501 11299 14535
rect 11241 14495 11299 14501
rect 11330 14492 11336 14544
rect 11388 14492 11394 14544
rect 13909 14535 13967 14541
rect 13909 14532 13921 14535
rect 11532 14504 12020 14532
rect 6273 14467 6331 14473
rect 6273 14433 6285 14467
rect 6319 14464 6331 14467
rect 6454 14464 6460 14476
rect 6319 14436 6460 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 9214 14424 9220 14476
rect 9272 14424 9278 14476
rect 9398 14424 9404 14476
rect 9456 14464 9462 14476
rect 9582 14464 9588 14476
rect 9456 14436 9588 14464
rect 9456 14424 9462 14436
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 9953 14467 10011 14473
rect 9953 14433 9965 14467
rect 9999 14464 10011 14467
rect 10042 14464 10048 14476
rect 9999 14436 10048 14464
rect 9999 14433 10011 14436
rect 9953 14427 10011 14433
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 10226 14424 10232 14476
rect 10284 14424 10290 14476
rect 10413 14467 10471 14473
rect 10413 14433 10425 14467
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 6362 14356 6368 14408
rect 6420 14396 6426 14408
rect 9030 14396 9036 14408
rect 6420 14368 9036 14396
rect 6420 14356 6426 14368
rect 9030 14356 9036 14368
rect 9088 14356 9094 14408
rect 9766 14356 9772 14408
rect 9824 14396 9830 14408
rect 10428 14396 10456 14427
rect 10870 14424 10876 14476
rect 10928 14464 10934 14476
rect 11532 14473 11560 14504
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 10928 14436 11161 14464
rect 10928 14424 10934 14436
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 11149 14427 11207 14433
rect 11517 14467 11575 14473
rect 11517 14433 11529 14467
rect 11563 14433 11575 14467
rect 11517 14427 11575 14433
rect 11606 14424 11612 14476
rect 11664 14464 11670 14476
rect 11992 14473 12020 14504
rect 13464 14504 13921 14532
rect 13464 14476 13492 14504
rect 13909 14501 13921 14504
rect 13955 14501 13967 14535
rect 14642 14532 14648 14544
rect 13909 14495 13967 14501
rect 14016 14504 14648 14532
rect 11885 14467 11943 14473
rect 11885 14464 11897 14467
rect 11664 14436 11897 14464
rect 11664 14424 11670 14436
rect 11885 14433 11897 14436
rect 11931 14433 11943 14467
rect 11885 14427 11943 14433
rect 11977 14467 12035 14473
rect 11977 14433 11989 14467
rect 12023 14464 12035 14467
rect 12342 14464 12348 14476
rect 12023 14436 12348 14464
rect 12023 14433 12035 14436
rect 11977 14427 12035 14433
rect 12342 14424 12348 14436
rect 12400 14424 12406 14476
rect 12805 14467 12863 14473
rect 12805 14433 12817 14467
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 9824 14368 10456 14396
rect 9824 14356 9830 14368
rect 11422 14356 11428 14408
rect 11480 14396 11486 14408
rect 11701 14399 11759 14405
rect 11701 14396 11713 14399
rect 11480 14368 11713 14396
rect 11480 14356 11486 14368
rect 11701 14365 11713 14368
rect 11747 14365 11759 14399
rect 12820 14396 12848 14427
rect 13078 14424 13084 14476
rect 13136 14424 13142 14476
rect 13357 14467 13415 14473
rect 13357 14433 13369 14467
rect 13403 14464 13415 14467
rect 13446 14464 13452 14476
rect 13403 14436 13452 14464
rect 13403 14433 13415 14436
rect 13357 14427 13415 14433
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 13817 14467 13875 14473
rect 13817 14464 13829 14467
rect 13587 14436 13829 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 13817 14433 13829 14436
rect 13863 14464 13875 14467
rect 14016 14464 14044 14504
rect 14642 14492 14648 14504
rect 14700 14492 14706 14544
rect 14844 14541 14872 14572
rect 15010 14560 15016 14612
rect 15068 14560 15074 14612
rect 17503 14603 17561 14609
rect 17503 14569 17515 14603
rect 17549 14600 17561 14603
rect 18690 14600 18696 14612
rect 17549 14572 18696 14600
rect 17549 14569 17561 14572
rect 17503 14563 17561 14569
rect 18690 14560 18696 14572
rect 18748 14560 18754 14612
rect 18874 14560 18880 14612
rect 18932 14600 18938 14612
rect 19061 14603 19119 14609
rect 19061 14600 19073 14603
rect 18932 14572 19073 14600
rect 18932 14560 18938 14572
rect 19061 14569 19073 14572
rect 19107 14569 19119 14603
rect 19061 14563 19119 14569
rect 21818 14560 21824 14612
rect 21876 14600 21882 14612
rect 22189 14603 22247 14609
rect 22189 14600 22201 14603
rect 21876 14572 22201 14600
rect 21876 14560 21882 14572
rect 22189 14569 22201 14572
rect 22235 14569 22247 14603
rect 22189 14563 22247 14569
rect 14737 14535 14795 14541
rect 14737 14501 14749 14535
rect 14783 14501 14795 14535
rect 14737 14495 14795 14501
rect 14829 14535 14887 14541
rect 14829 14501 14841 14535
rect 14875 14501 14887 14535
rect 14829 14495 14887 14501
rect 13863 14436 14044 14464
rect 13863 14433 13875 14436
rect 13817 14427 13875 14433
rect 11701 14359 11759 14365
rect 12406 14368 12848 14396
rect 13265 14399 13323 14405
rect 12406 14340 12434 14368
rect 13265 14365 13277 14399
rect 13311 14396 13323 14399
rect 13556 14396 13584 14427
rect 14090 14424 14096 14476
rect 14148 14424 14154 14476
rect 14752 14464 14780 14495
rect 15028 14464 15056 14560
rect 17586 14492 17592 14544
rect 17644 14492 17650 14544
rect 19213 14535 19271 14541
rect 19213 14532 19225 14535
rect 17696 14504 19225 14532
rect 17696 14476 17724 14504
rect 19213 14501 19225 14504
rect 19259 14501 19271 14535
rect 19213 14495 19271 14501
rect 19429 14535 19487 14541
rect 19429 14501 19441 14535
rect 19475 14501 19487 14535
rect 19429 14495 19487 14501
rect 14752 14436 15056 14464
rect 15105 14467 15163 14473
rect 15105 14433 15117 14467
rect 15151 14433 15163 14467
rect 15105 14427 15163 14433
rect 15120 14396 15148 14427
rect 16574 14424 16580 14476
rect 16632 14464 16638 14476
rect 16669 14467 16727 14473
rect 16669 14464 16681 14467
rect 16632 14436 16681 14464
rect 16632 14424 16638 14436
rect 16669 14433 16681 14436
rect 16715 14433 16727 14467
rect 16669 14427 16727 14433
rect 17402 14424 17408 14476
rect 17460 14424 17466 14476
rect 17678 14424 17684 14476
rect 17736 14424 17742 14476
rect 17773 14467 17831 14473
rect 17773 14433 17785 14467
rect 17819 14433 17831 14467
rect 17773 14427 17831 14433
rect 13311 14368 13584 14396
rect 14568 14368 15148 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 9401 14331 9459 14337
rect 9401 14297 9413 14331
rect 9447 14328 9459 14331
rect 10226 14328 10232 14340
rect 9447 14300 10232 14328
rect 9447 14297 9459 14300
rect 9401 14291 9459 14297
rect 10226 14288 10232 14300
rect 10284 14288 10290 14340
rect 10965 14331 11023 14337
rect 10965 14297 10977 14331
rect 11011 14328 11023 14331
rect 12342 14328 12348 14340
rect 11011 14300 12348 14328
rect 11011 14297 11023 14300
rect 10965 14291 11023 14297
rect 12342 14288 12348 14300
rect 12400 14300 12434 14340
rect 14568 14328 14596 14368
rect 16942 14356 16948 14408
rect 17000 14396 17006 14408
rect 17494 14396 17500 14408
rect 17000 14368 17500 14396
rect 17000 14356 17006 14368
rect 17494 14356 17500 14368
rect 17552 14356 17558 14408
rect 17788 14396 17816 14427
rect 17954 14424 17960 14476
rect 18012 14424 18018 14476
rect 18598 14424 18604 14476
rect 18656 14424 18662 14476
rect 18046 14396 18052 14408
rect 17788 14368 18052 14396
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 18138 14356 18144 14408
rect 18196 14356 18202 14408
rect 18414 14356 18420 14408
rect 18472 14396 18478 14408
rect 18509 14399 18567 14405
rect 18509 14396 18521 14399
rect 18472 14368 18521 14396
rect 18472 14356 18478 14368
rect 18509 14365 18521 14368
rect 18555 14365 18567 14399
rect 19444 14396 19472 14495
rect 22094 14492 22100 14544
rect 22152 14532 22158 14544
rect 22557 14535 22615 14541
rect 22557 14532 22569 14535
rect 22152 14504 22569 14532
rect 22152 14492 22158 14504
rect 22557 14501 22569 14504
rect 22603 14501 22615 14535
rect 22557 14495 22615 14501
rect 22649 14535 22707 14541
rect 22649 14501 22661 14535
rect 22695 14532 22707 14535
rect 22922 14532 22928 14544
rect 22695 14504 22928 14532
rect 22695 14501 22707 14504
rect 22649 14495 22707 14501
rect 22922 14492 22928 14504
rect 22980 14492 22986 14544
rect 21542 14424 21548 14476
rect 21600 14424 21606 14476
rect 22005 14467 22063 14473
rect 22005 14433 22017 14467
rect 22051 14464 22063 14467
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 22051 14436 22293 14464
rect 22051 14433 22063 14436
rect 22005 14427 22063 14433
rect 22281 14433 22293 14436
rect 22327 14433 22339 14467
rect 22281 14427 22339 14433
rect 22370 14424 22376 14476
rect 22428 14464 22434 14476
rect 22465 14467 22523 14473
rect 22465 14464 22477 14467
rect 22428 14436 22477 14464
rect 22428 14424 22434 14436
rect 22465 14433 22477 14436
rect 22511 14433 22523 14467
rect 22465 14427 22523 14433
rect 22738 14424 22744 14476
rect 22796 14473 22802 14476
rect 22796 14467 22825 14473
rect 22813 14433 22825 14467
rect 22796 14427 22825 14433
rect 22796 14424 22802 14427
rect 18509 14359 18567 14365
rect 18800 14368 19472 14396
rect 14292 14300 14596 14328
rect 12400 14288 12406 14300
rect 14292 14272 14320 14300
rect 5813 14263 5871 14269
rect 5813 14229 5825 14263
rect 5859 14260 5871 14263
rect 5994 14260 6000 14272
rect 5859 14232 6000 14260
rect 5859 14229 5871 14232
rect 5813 14223 5871 14229
rect 5994 14220 6000 14232
rect 6052 14220 6058 14272
rect 9493 14263 9551 14269
rect 9493 14229 9505 14263
rect 9539 14260 9551 14263
rect 9950 14260 9956 14272
rect 9539 14232 9956 14260
rect 9539 14229 9551 14232
rect 9493 14223 9551 14229
rect 9950 14220 9956 14232
rect 10008 14220 10014 14272
rect 10134 14220 10140 14272
rect 10192 14260 10198 14272
rect 10870 14260 10876 14272
rect 10192 14232 10876 14260
rect 10192 14220 10198 14232
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 11790 14220 11796 14272
rect 11848 14220 11854 14272
rect 13449 14263 13507 14269
rect 13449 14229 13461 14263
rect 13495 14260 13507 14263
rect 13722 14260 13728 14272
rect 13495 14232 13728 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 14274 14220 14280 14272
rect 14332 14220 14338 14272
rect 14366 14220 14372 14272
rect 14424 14220 14430 14272
rect 14568 14269 14596 14300
rect 16853 14331 16911 14337
rect 16853 14297 16865 14331
rect 16899 14328 16911 14331
rect 18322 14328 18328 14340
rect 16899 14300 18328 14328
rect 16899 14297 16911 14300
rect 16853 14291 16911 14297
rect 18322 14288 18328 14300
rect 18380 14288 18386 14340
rect 14553 14263 14611 14269
rect 14553 14229 14565 14263
rect 14599 14229 14611 14263
rect 14553 14223 14611 14229
rect 14642 14220 14648 14272
rect 14700 14260 14706 14272
rect 14829 14263 14887 14269
rect 14829 14260 14841 14263
rect 14700 14232 14841 14260
rect 14700 14220 14706 14232
rect 14829 14229 14841 14232
rect 14875 14229 14887 14263
rect 14829 14223 14887 14229
rect 16758 14220 16764 14272
rect 16816 14220 16822 14272
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 18800 14260 18828 14368
rect 21910 14356 21916 14408
rect 21968 14356 21974 14408
rect 22925 14399 22983 14405
rect 22925 14365 22937 14399
rect 22971 14365 22983 14399
rect 22925 14359 22983 14365
rect 22462 14328 22468 14340
rect 22020 14300 22468 14328
rect 17460 14232 18828 14260
rect 18877 14263 18935 14269
rect 17460 14220 17466 14232
rect 18877 14229 18889 14263
rect 18923 14260 18935 14263
rect 18966 14260 18972 14272
rect 18923 14232 18972 14260
rect 18923 14229 18935 14232
rect 18877 14223 18935 14229
rect 18966 14220 18972 14232
rect 19024 14220 19030 14272
rect 19242 14220 19248 14272
rect 19300 14220 19306 14272
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 20806 14260 20812 14272
rect 19392 14232 20812 14260
rect 19392 14220 19398 14232
rect 20806 14220 20812 14232
rect 20864 14220 20870 14272
rect 22020 14269 22048 14300
rect 22462 14288 22468 14300
rect 22520 14288 22526 14340
rect 22830 14288 22836 14340
rect 22888 14328 22894 14340
rect 22940 14328 22968 14359
rect 22888 14300 22968 14328
rect 22888 14288 22894 14300
rect 22005 14263 22063 14269
rect 22005 14229 22017 14263
rect 22051 14229 22063 14263
rect 22005 14223 22063 14229
rect 552 14170 23368 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 23368 14170
rect 552 14096 23368 14118
rect 4249 14059 4307 14065
rect 4249 14025 4261 14059
rect 4295 14056 4307 14059
rect 6178 14056 6184 14068
rect 4295 14028 6184 14056
rect 4295 14025 4307 14028
rect 4249 14019 4307 14025
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 8941 14059 8999 14065
rect 8941 14025 8953 14059
rect 8987 14056 8999 14059
rect 9582 14056 9588 14068
rect 8987 14028 9588 14056
rect 8987 14025 8999 14028
rect 8941 14019 8999 14025
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 10965 14059 11023 14065
rect 10965 14025 10977 14059
rect 11011 14056 11023 14059
rect 11330 14056 11336 14068
rect 11011 14028 11336 14056
rect 11011 14025 11023 14028
rect 10965 14019 11023 14025
rect 5721 13991 5779 13997
rect 5721 13957 5733 13991
rect 5767 13957 5779 13991
rect 5721 13951 5779 13957
rect 7193 13991 7251 13997
rect 7193 13957 7205 13991
rect 7239 13957 7251 13991
rect 7193 13951 7251 13957
rect 5373 13855 5431 13861
rect 5373 13821 5385 13855
rect 5419 13852 5431 13855
rect 5534 13852 5540 13864
rect 5419 13824 5540 13852
rect 5419 13821 5431 13824
rect 5373 13815 5431 13821
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 5629 13855 5687 13861
rect 5629 13821 5641 13855
rect 5675 13821 5687 13855
rect 5736 13852 5764 13951
rect 7208 13920 7236 13951
rect 9214 13948 9220 14000
rect 9272 13948 9278 14000
rect 10042 13948 10048 14000
rect 10100 13988 10106 14000
rect 10100 13960 10732 13988
rect 10100 13948 10106 13960
rect 7024 13892 7236 13920
rect 6845 13855 6903 13861
rect 5736 13824 6776 13852
rect 5629 13815 5687 13821
rect 5644 13716 5672 13815
rect 6748 13784 6776 13824
rect 6845 13821 6857 13855
rect 6891 13852 6903 13855
rect 7024 13852 7052 13892
rect 7650 13880 7656 13932
rect 7708 13880 7714 13932
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 8110 13920 8116 13932
rect 7883 13892 8116 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 9232 13920 9260 13948
rect 9140 13892 9260 13920
rect 9784 13892 10272 13920
rect 6891 13824 7052 13852
rect 6891 13821 6903 13824
rect 6845 13815 6903 13821
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 8941 13855 8999 13861
rect 7156 13824 7696 13852
rect 7156 13812 7162 13824
rect 7006 13784 7012 13796
rect 6748 13756 7012 13784
rect 7006 13744 7012 13756
rect 7064 13784 7070 13796
rect 7561 13787 7619 13793
rect 7561 13784 7573 13787
rect 7064 13756 7573 13784
rect 7064 13744 7070 13756
rect 7561 13753 7573 13756
rect 7607 13753 7619 13787
rect 7561 13747 7619 13753
rect 5810 13716 5816 13728
rect 5644 13688 5816 13716
rect 5810 13676 5816 13688
rect 5868 13716 5874 13728
rect 7098 13716 7104 13728
rect 5868 13688 7104 13716
rect 5868 13676 5874 13688
rect 7098 13676 7104 13688
rect 7156 13676 7162 13728
rect 7668 13716 7696 13824
rect 8941 13821 8953 13855
rect 8987 13852 8999 13855
rect 9030 13852 9036 13864
rect 8987 13824 9036 13852
rect 8987 13821 8999 13824
rect 8941 13815 8999 13821
rect 9030 13812 9036 13824
rect 9088 13812 9094 13864
rect 9140 13861 9168 13892
rect 9784 13864 9812 13892
rect 9125 13855 9183 13861
rect 9125 13821 9137 13855
rect 9171 13821 9183 13855
rect 9125 13815 9183 13821
rect 9217 13855 9275 13861
rect 9217 13821 9229 13855
rect 9263 13852 9275 13855
rect 9398 13852 9404 13864
rect 9263 13824 9404 13852
rect 9263 13821 9275 13824
rect 9217 13815 9275 13821
rect 9398 13812 9404 13824
rect 9456 13812 9462 13864
rect 9766 13812 9772 13864
rect 9824 13812 9830 13864
rect 9950 13812 9956 13864
rect 10008 13852 10014 13864
rect 10244 13861 10272 13892
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 10008 13824 10057 13852
rect 10008 13812 10014 13824
rect 10045 13821 10057 13824
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 10229 13855 10287 13861
rect 10229 13821 10241 13855
rect 10275 13821 10287 13855
rect 10229 13815 10287 13821
rect 10594 13812 10600 13864
rect 10652 13812 10658 13864
rect 10704 13852 10732 13960
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13920 10839 13923
rect 10980 13920 11008 14019
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 14642 14016 14648 14068
rect 14700 14016 14706 14068
rect 16942 14016 16948 14068
rect 17000 14016 17006 14068
rect 17313 14059 17371 14065
rect 17313 14025 17325 14059
rect 17359 14056 17371 14059
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17359 14028 17785 14056
rect 17359 14025 17371 14028
rect 17313 14019 17371 14025
rect 17773 14025 17785 14028
rect 17819 14056 17831 14059
rect 17862 14056 17868 14068
rect 17819 14028 17868 14056
rect 17819 14025 17831 14028
rect 17773 14019 17831 14025
rect 17862 14016 17868 14028
rect 17920 14016 17926 14068
rect 17954 14016 17960 14068
rect 18012 14016 18018 14068
rect 18046 14016 18052 14068
rect 18104 14016 18110 14068
rect 19058 14016 19064 14068
rect 19116 14016 19122 14068
rect 19245 14059 19303 14065
rect 19245 14025 19257 14059
rect 19291 14056 19303 14059
rect 20530 14056 20536 14068
rect 19291 14028 20536 14056
rect 19291 14025 19303 14028
rect 19245 14019 19303 14025
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 21450 14016 21456 14068
rect 21508 14056 21514 14068
rect 21729 14059 21787 14065
rect 21729 14056 21741 14059
rect 21508 14028 21741 14056
rect 21508 14016 21514 14028
rect 21729 14025 21741 14028
rect 21775 14025 21787 14059
rect 21729 14019 21787 14025
rect 21910 14016 21916 14068
rect 21968 14016 21974 14068
rect 13814 13948 13820 14000
rect 13872 13988 13878 14000
rect 14737 13991 14795 13997
rect 14737 13988 14749 13991
rect 13872 13960 14749 13988
rect 13872 13948 13878 13960
rect 14737 13957 14749 13960
rect 14783 13957 14795 13991
rect 19334 13988 19340 14000
rect 14737 13951 14795 13957
rect 16500 13960 19340 13988
rect 10827 13892 11008 13920
rect 10827 13889 10839 13892
rect 10781 13883 10839 13889
rect 12342 13880 12348 13932
rect 12400 13920 12406 13932
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 12400 13892 13093 13920
rect 12400 13880 12406 13892
rect 13081 13889 13093 13892
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13170 13880 13176 13932
rect 13228 13880 13234 13932
rect 13262 13880 13268 13932
rect 13320 13920 13326 13932
rect 14829 13923 14887 13929
rect 13320 13892 14780 13920
rect 13320 13880 13326 13892
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10704 13824 10885 13852
rect 10873 13821 10885 13824
rect 10919 13821 10931 13855
rect 10873 13815 10931 13821
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11057 13855 11115 13861
rect 11057 13852 11069 13855
rect 11020 13824 11069 13852
rect 11020 13812 11026 13824
rect 11057 13821 11069 13824
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 12986 13812 12992 13864
rect 13044 13812 13050 13864
rect 13722 13812 13728 13864
rect 13780 13812 13786 13864
rect 13879 13855 13937 13861
rect 13879 13821 13891 13855
rect 13925 13852 13937 13855
rect 14090 13852 14096 13864
rect 13925 13824 14096 13852
rect 13925 13821 13937 13824
rect 13879 13815 13937 13821
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 14553 13855 14611 13861
rect 14553 13852 14565 13855
rect 14424 13824 14565 13852
rect 14424 13812 14430 13824
rect 14553 13821 14565 13824
rect 14599 13821 14611 13855
rect 14752 13852 14780 13892
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 14918 13920 14924 13932
rect 14875 13892 14924 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 15396 13892 15608 13920
rect 15396 13852 15424 13892
rect 14752 13824 15424 13852
rect 14553 13815 14611 13821
rect 15470 13812 15476 13864
rect 15528 13812 15534 13864
rect 15580 13852 15608 13892
rect 16500 13852 16528 13960
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 18138 13880 18144 13932
rect 18196 13920 18202 13932
rect 18877 13923 18935 13929
rect 18877 13920 18889 13923
rect 18196 13892 18889 13920
rect 18196 13880 18202 13892
rect 18877 13889 18889 13892
rect 18923 13889 18935 13923
rect 18877 13883 18935 13889
rect 19978 13880 19984 13932
rect 20036 13920 20042 13932
rect 20349 13923 20407 13929
rect 20349 13920 20361 13923
rect 20036 13892 20361 13920
rect 20036 13880 20042 13892
rect 20349 13889 20361 13892
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 15580 13824 16528 13852
rect 16758 13812 16764 13864
rect 16816 13852 16822 13864
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 16816 13824 16957 13852
rect 16816 13812 16822 13824
rect 16945 13821 16957 13824
rect 16991 13821 17003 13855
rect 16945 13815 17003 13821
rect 17037 13855 17095 13861
rect 17037 13821 17049 13855
rect 17083 13821 17095 13855
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17037 13815 17095 13821
rect 17604 13824 18061 13852
rect 13078 13784 13084 13796
rect 9048 13756 13084 13784
rect 9048 13716 9076 13756
rect 13078 13744 13084 13756
rect 13136 13744 13142 13796
rect 15740 13787 15798 13793
rect 15740 13753 15752 13787
rect 15786 13784 15798 13787
rect 16114 13784 16120 13796
rect 15786 13756 16120 13784
rect 15786 13753 15798 13756
rect 15740 13747 15798 13753
rect 16114 13744 16120 13756
rect 16172 13744 16178 13796
rect 17052 13784 17080 13815
rect 17604 13796 17632 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18322 13852 18328 13864
rect 18049 13815 18107 13821
rect 18156 13824 18328 13852
rect 16868 13756 17080 13784
rect 7668 13688 9076 13716
rect 9490 13676 9496 13728
rect 9548 13716 9554 13728
rect 9585 13719 9643 13725
rect 9585 13716 9597 13719
rect 9548 13688 9597 13716
rect 9548 13676 9554 13688
rect 9585 13685 9597 13688
rect 9631 13685 9643 13719
rect 9585 13679 9643 13685
rect 10134 13676 10140 13728
rect 10192 13676 10198 13728
rect 10410 13676 10416 13728
rect 10468 13676 10474 13728
rect 12802 13676 12808 13728
rect 12860 13676 12866 13728
rect 14090 13676 14096 13728
rect 14148 13676 14154 13728
rect 16574 13676 16580 13728
rect 16632 13716 16638 13728
rect 16868 13725 16896 13756
rect 17586 13744 17592 13796
rect 17644 13744 17650 13796
rect 17805 13787 17863 13793
rect 17805 13753 17817 13787
rect 17851 13784 17863 13787
rect 18156 13784 18184 13824
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 18782 13812 18788 13864
rect 18840 13812 18846 13864
rect 18966 13812 18972 13864
rect 19024 13852 19030 13864
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 19024 13824 19073 13852
rect 19024 13812 19030 13824
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 19886 13812 19892 13864
rect 19944 13852 19950 13864
rect 20073 13855 20131 13861
rect 20073 13852 20085 13855
rect 19944 13824 20085 13852
rect 19944 13812 19950 13824
rect 20073 13821 20085 13824
rect 20119 13821 20131 13855
rect 20073 13815 20131 13821
rect 17851 13756 18184 13784
rect 17851 13753 17863 13756
rect 17805 13747 17863 13753
rect 16853 13719 16911 13725
rect 16853 13716 16865 13719
rect 16632 13688 16865 13716
rect 16632 13676 16638 13688
rect 16853 13685 16865 13688
rect 16899 13685 16911 13719
rect 16853 13679 16911 13685
rect 17954 13676 17960 13728
rect 18012 13716 18018 13728
rect 18233 13719 18291 13725
rect 18233 13716 18245 13719
rect 18012 13688 18245 13716
rect 18012 13676 18018 13688
rect 18233 13685 18245 13688
rect 18279 13685 18291 13719
rect 18233 13679 18291 13685
rect 19886 13676 19892 13728
rect 19944 13676 19950 13728
rect 20088 13716 20116 13815
rect 20254 13812 20260 13864
rect 20312 13812 20318 13864
rect 20616 13855 20674 13861
rect 20616 13821 20628 13855
rect 20662 13852 20674 13855
rect 21082 13852 21088 13864
rect 20662 13824 21088 13852
rect 20662 13821 20674 13824
rect 20616 13815 20674 13821
rect 21082 13812 21088 13824
rect 21140 13812 21146 13864
rect 22094 13812 22100 13864
rect 22152 13812 22158 13864
rect 22189 13855 22247 13861
rect 22189 13821 22201 13855
rect 22235 13852 22247 13855
rect 22278 13852 22284 13864
rect 22235 13824 22284 13852
rect 22235 13821 22247 13824
rect 22189 13815 22247 13821
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 21913 13787 21971 13793
rect 21913 13753 21925 13787
rect 21959 13784 21971 13787
rect 21959 13756 22140 13784
rect 21959 13753 21971 13756
rect 21913 13747 21971 13753
rect 22112 13728 22140 13756
rect 20530 13716 20536 13728
rect 20088 13688 20536 13716
rect 20530 13676 20536 13688
rect 20588 13676 20594 13728
rect 22094 13676 22100 13728
rect 22152 13676 22158 13728
rect 552 13626 23368 13648
rect 552 13574 4322 13626
rect 4374 13574 4386 13626
rect 4438 13574 4450 13626
rect 4502 13574 4514 13626
rect 4566 13574 4578 13626
rect 4630 13574 23368 13626
rect 552 13552 23368 13574
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 5592 13484 5825 13512
rect 5592 13472 5598 13484
rect 5813 13481 5825 13484
rect 5859 13481 5871 13515
rect 5813 13475 5871 13481
rect 6178 13472 6184 13524
rect 6236 13472 6242 13524
rect 10134 13512 10140 13524
rect 8772 13484 10140 13512
rect 5718 13404 5724 13456
rect 5776 13444 5782 13456
rect 6273 13447 6331 13453
rect 6273 13444 6285 13447
rect 5776 13416 6285 13444
rect 5776 13404 5782 13416
rect 6273 13413 6285 13416
rect 6319 13413 6331 13447
rect 8110 13444 8116 13456
rect 6273 13407 6331 13413
rect 6472 13416 8116 13444
rect 6472 13317 6500 13416
rect 8110 13404 8116 13416
rect 8168 13404 8174 13456
rect 7009 13379 7067 13385
rect 7009 13345 7021 13379
rect 7055 13376 7067 13379
rect 7098 13376 7104 13388
rect 7055 13348 7104 13376
rect 7055 13345 7067 13348
rect 7009 13339 7067 13345
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 7282 13385 7288 13388
rect 7276 13339 7288 13385
rect 7282 13336 7288 13339
rect 7340 13336 7346 13388
rect 8772 13385 8800 13484
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 12342 13512 12348 13524
rect 11900 13484 12348 13512
rect 9490 13444 9496 13456
rect 8956 13416 9496 13444
rect 8956 13385 8984 13416
rect 9490 13404 9496 13416
rect 9548 13444 9554 13456
rect 9548 13416 9996 13444
rect 9548 13404 9554 13416
rect 8757 13379 8815 13385
rect 8757 13345 8769 13379
rect 8803 13345 8815 13379
rect 8757 13339 8815 13345
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 9214 13336 9220 13388
rect 9272 13336 9278 13388
rect 9306 13336 9312 13388
rect 9364 13336 9370 13388
rect 9401 13379 9459 13385
rect 9401 13345 9413 13379
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 9416 13308 9444 13339
rect 9582 13336 9588 13388
rect 9640 13336 9646 13388
rect 9968 13385 9996 13416
rect 9953 13379 10011 13385
rect 9953 13345 9965 13379
rect 9999 13345 10011 13379
rect 9953 13339 10011 13345
rect 10226 13336 10232 13388
rect 10284 13336 10290 13388
rect 11790 13336 11796 13388
rect 11848 13336 11854 13388
rect 11900 13385 11928 13484
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 13262 13512 13268 13524
rect 12492 13484 13268 13512
rect 12492 13472 12498 13484
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 16114 13472 16120 13524
rect 16172 13472 16178 13524
rect 18138 13472 18144 13524
rect 18196 13512 18202 13524
rect 18525 13515 18583 13521
rect 18525 13512 18537 13515
rect 18196 13484 18537 13512
rect 18196 13472 18202 13484
rect 18525 13481 18537 13484
rect 18571 13481 18583 13515
rect 18525 13475 18583 13481
rect 21744 13484 22094 13512
rect 16485 13447 16543 13453
rect 11992 13416 16436 13444
rect 11885 13379 11943 13385
rect 11885 13345 11897 13379
rect 11931 13345 11943 13379
rect 11885 13339 11943 13345
rect 11992 13320 12020 13416
rect 12345 13379 12403 13385
rect 12345 13345 12357 13379
rect 12391 13345 12403 13379
rect 12345 13339 12403 13345
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9416 13280 9689 13308
rect 6457 13271 6515 13277
rect 9677 13277 9689 13280
rect 9723 13308 9735 13311
rect 10321 13311 10379 13317
rect 10321 13308 10333 13311
rect 9723 13280 10333 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 10321 13277 10333 13280
rect 10367 13277 10379 13311
rect 10321 13271 10379 13277
rect 11974 13268 11980 13320
rect 12032 13268 12038 13320
rect 12066 13268 12072 13320
rect 12124 13268 12130 13320
rect 12360 13308 12388 13339
rect 12802 13336 12808 13388
rect 12860 13336 12866 13388
rect 12897 13379 12955 13385
rect 12897 13345 12909 13379
rect 12943 13376 12955 13379
rect 13722 13376 13728 13388
rect 12943 13348 13728 13376
rect 12943 13345 12955 13348
rect 12897 13339 12955 13345
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 14090 13336 14096 13388
rect 14148 13376 14154 13388
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 14148 13348 14289 13376
rect 14148 13336 14154 13348
rect 14277 13345 14289 13348
rect 14323 13345 14335 13379
rect 14277 13339 14335 13345
rect 14366 13336 14372 13388
rect 14424 13336 14430 13388
rect 14461 13379 14519 13385
rect 14461 13345 14473 13379
rect 14507 13376 14519 13379
rect 14826 13376 14832 13388
rect 14507 13348 14832 13376
rect 14507 13345 14519 13348
rect 14461 13339 14519 13345
rect 12526 13308 12532 13320
rect 12360 13280 12532 13308
rect 12526 13268 12532 13280
rect 12584 13268 12590 13320
rect 13906 13268 13912 13320
rect 13964 13308 13970 13320
rect 14476 13308 14504 13339
rect 14826 13336 14832 13348
rect 14884 13336 14890 13388
rect 14921 13379 14979 13385
rect 14921 13345 14933 13379
rect 14967 13345 14979 13379
rect 16408 13376 16436 13416
rect 16485 13413 16497 13447
rect 16531 13444 16543 13447
rect 16574 13444 16580 13456
rect 16531 13416 16580 13444
rect 16531 13413 16543 13416
rect 16485 13407 16543 13413
rect 16574 13404 16580 13416
rect 16632 13404 16638 13456
rect 17402 13404 17408 13456
rect 17460 13444 17466 13456
rect 17862 13444 17868 13456
rect 17460 13416 17868 13444
rect 17460 13404 17466 13416
rect 17862 13404 17868 13416
rect 17920 13444 17926 13456
rect 18325 13447 18383 13453
rect 18325 13444 18337 13447
rect 17920 13416 18337 13444
rect 17920 13404 17926 13416
rect 18325 13413 18337 13416
rect 18371 13413 18383 13447
rect 18325 13407 18383 13413
rect 19242 13404 19248 13456
rect 19300 13444 19306 13456
rect 19889 13447 19947 13453
rect 19889 13444 19901 13447
rect 19300 13416 19901 13444
rect 19300 13404 19306 13416
rect 19889 13413 19901 13416
rect 19935 13413 19947 13447
rect 19889 13407 19947 13413
rect 20714 13404 20720 13456
rect 20772 13404 20778 13456
rect 20898 13404 20904 13456
rect 20956 13444 20962 13456
rect 21174 13444 21180 13456
rect 20956 13416 21180 13444
rect 20956 13404 20962 13416
rect 21174 13404 21180 13416
rect 21232 13444 21238 13456
rect 21744 13453 21772 13484
rect 22066 13456 22094 13484
rect 21269 13447 21327 13453
rect 21269 13444 21281 13447
rect 21232 13416 21281 13444
rect 21232 13404 21238 13416
rect 21269 13413 21281 13416
rect 21315 13413 21327 13447
rect 21469 13447 21527 13453
rect 21469 13444 21481 13447
rect 21269 13407 21327 13413
rect 21376 13416 21481 13444
rect 20162 13376 20168 13388
rect 16408 13348 20168 13376
rect 14921 13339 14979 13345
rect 13964 13280 14504 13308
rect 14553 13311 14611 13317
rect 13964 13268 13970 13280
rect 14553 13277 14565 13311
rect 14599 13308 14611 13311
rect 14737 13311 14795 13317
rect 14737 13308 14749 13311
rect 14599 13280 14749 13308
rect 14599 13277 14611 13280
rect 14553 13271 14611 13277
rect 14737 13277 14749 13280
rect 14783 13277 14795 13311
rect 14737 13271 14795 13277
rect 8849 13243 8907 13249
rect 8849 13209 8861 13243
rect 8895 13240 8907 13243
rect 9306 13240 9312 13252
rect 8895 13212 9312 13240
rect 8895 13209 8907 13212
rect 8849 13203 8907 13209
rect 9306 13200 9312 13212
rect 9364 13240 9370 13252
rect 9769 13243 9827 13249
rect 9769 13240 9781 13243
rect 9364 13212 9781 13240
rect 9364 13200 9370 13212
rect 9769 13209 9781 13212
rect 9815 13209 9827 13243
rect 14936 13240 14964 13339
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 20257 13379 20315 13385
rect 20257 13345 20269 13379
rect 20303 13376 20315 13379
rect 20732 13376 20760 13404
rect 21376 13376 21404 13416
rect 21469 13413 21481 13416
rect 21515 13413 21527 13447
rect 21469 13407 21527 13413
rect 21729 13447 21787 13453
rect 21729 13413 21741 13447
rect 21775 13413 21787 13447
rect 21929 13447 21987 13453
rect 21929 13444 21941 13447
rect 21729 13407 21787 13413
rect 21836 13416 21941 13444
rect 20303 13348 21404 13376
rect 20303 13345 20315 13348
rect 20257 13339 20315 13345
rect 21634 13336 21640 13388
rect 21692 13376 21698 13388
rect 21836 13376 21864 13416
rect 21929 13413 21941 13416
rect 21975 13413 21987 13447
rect 22066 13416 22100 13456
rect 21929 13407 21987 13413
rect 22094 13404 22100 13416
rect 22152 13444 22158 13456
rect 22922 13444 22928 13456
rect 22152 13416 22928 13444
rect 22152 13404 22158 13416
rect 22922 13404 22928 13416
rect 22980 13404 22986 13456
rect 22373 13379 22431 13385
rect 22373 13376 22385 13379
rect 21692 13348 21864 13376
rect 22066 13348 22385 13376
rect 21692 13336 21698 13348
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13308 15163 13311
rect 15286 13308 15292 13320
rect 15151 13280 15292 13308
rect 15151 13277 15163 13280
rect 15105 13271 15163 13277
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 16390 13268 16396 13320
rect 16448 13308 16454 13320
rect 16577 13311 16635 13317
rect 16577 13308 16589 13311
rect 16448 13280 16589 13308
rect 16448 13268 16454 13280
rect 16577 13277 16589 13280
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 16761 13311 16819 13317
rect 16761 13277 16773 13311
rect 16807 13308 16819 13311
rect 16850 13308 16856 13320
rect 16807 13280 16856 13308
rect 16807 13277 16819 13280
rect 16761 13271 16819 13277
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 20441 13311 20499 13317
rect 20441 13277 20453 13311
rect 20487 13277 20499 13311
rect 20441 13271 20499 13277
rect 16482 13240 16488 13252
rect 14936 13212 16488 13240
rect 9769 13203 9827 13209
rect 16482 13200 16488 13212
rect 16540 13200 16546 13252
rect 18693 13243 18751 13249
rect 18693 13209 18705 13243
rect 18739 13240 18751 13243
rect 19334 13240 19340 13252
rect 18739 13212 19340 13240
rect 18739 13209 18751 13212
rect 18693 13203 18751 13209
rect 19334 13200 19340 13212
rect 19392 13240 19398 13252
rect 20456 13240 20484 13271
rect 20530 13268 20536 13320
rect 20588 13268 20594 13320
rect 20622 13268 20628 13320
rect 20680 13268 20686 13320
rect 20717 13311 20775 13317
rect 20717 13277 20729 13311
rect 20763 13308 20775 13311
rect 20806 13308 20812 13320
rect 20763 13280 20812 13308
rect 20763 13277 20775 13280
rect 20717 13271 20775 13277
rect 20806 13268 20812 13280
rect 20864 13268 20870 13320
rect 21818 13268 21824 13320
rect 21876 13308 21882 13320
rect 22066 13308 22094 13348
rect 22373 13345 22385 13348
rect 22419 13345 22431 13379
rect 22373 13339 22431 13345
rect 22557 13379 22615 13385
rect 22557 13345 22569 13379
rect 22603 13376 22615 13379
rect 22833 13379 22891 13385
rect 22833 13376 22845 13379
rect 22603 13348 22845 13376
rect 22603 13345 22615 13348
rect 22557 13339 22615 13345
rect 22833 13345 22845 13348
rect 22879 13345 22891 13379
rect 22833 13339 22891 13345
rect 21876 13280 22094 13308
rect 21876 13268 21882 13280
rect 22186 13268 22192 13320
rect 22244 13268 22250 13320
rect 22370 13240 22376 13252
rect 19392 13212 20300 13240
rect 20456 13212 21496 13240
rect 19392 13200 19398 13212
rect 20272 13184 20300 13212
rect 21468 13184 21496 13212
rect 21928 13212 22376 13240
rect 8386 13132 8392 13184
rect 8444 13132 8450 13184
rect 9030 13132 9036 13184
rect 9088 13132 9094 13184
rect 10134 13132 10140 13184
rect 10192 13132 10198 13184
rect 11606 13132 11612 13184
rect 11664 13132 11670 13184
rect 12710 13132 12716 13184
rect 12768 13132 12774 13184
rect 14093 13175 14151 13181
rect 14093 13141 14105 13175
rect 14139 13172 14151 13175
rect 14182 13172 14188 13184
rect 14139 13144 14188 13172
rect 14139 13141 14151 13144
rect 14093 13135 14151 13141
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 18509 13175 18567 13181
rect 18509 13141 18521 13175
rect 18555 13172 18567 13175
rect 18598 13172 18604 13184
rect 18555 13144 18604 13172
rect 18555 13141 18567 13144
rect 18509 13135 18567 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 19702 13132 19708 13184
rect 19760 13132 19766 13184
rect 19886 13132 19892 13184
rect 19944 13132 19950 13184
rect 20254 13132 20260 13184
rect 20312 13172 20318 13184
rect 20806 13172 20812 13184
rect 20312 13144 20812 13172
rect 20312 13132 20318 13144
rect 20806 13132 20812 13144
rect 20864 13132 20870 13184
rect 20901 13175 20959 13181
rect 20901 13141 20913 13175
rect 20947 13172 20959 13175
rect 21266 13172 21272 13184
rect 20947 13144 21272 13172
rect 20947 13141 20959 13144
rect 20901 13135 20959 13141
rect 21266 13132 21272 13144
rect 21324 13132 21330 13184
rect 21450 13132 21456 13184
rect 21508 13132 21514 13184
rect 21634 13132 21640 13184
rect 21692 13132 21698 13184
rect 21928 13181 21956 13212
rect 22370 13200 22376 13212
rect 22428 13200 22434 13252
rect 22646 13200 22652 13252
rect 22704 13200 22710 13252
rect 21913 13175 21971 13181
rect 21913 13141 21925 13175
rect 21959 13141 21971 13175
rect 21913 13135 21971 13141
rect 22094 13132 22100 13184
rect 22152 13132 22158 13184
rect 552 13082 23368 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 23368 13082
rect 552 13008 23368 13030
rect 6362 12928 6368 12980
rect 6420 12968 6426 12980
rect 6546 12968 6552 12980
rect 6420 12940 6552 12968
rect 6420 12928 6426 12940
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 7282 12928 7288 12980
rect 7340 12968 7346 12980
rect 7469 12971 7527 12977
rect 7469 12968 7481 12971
rect 7340 12940 7481 12968
rect 7340 12928 7346 12940
rect 7469 12937 7481 12940
rect 7515 12937 7527 12971
rect 11054 12968 11060 12980
rect 7469 12931 7527 12937
rect 8312 12940 11060 12968
rect 7098 12900 7104 12912
rect 6288 12872 7104 12900
rect 6288 12841 6316 12872
rect 7098 12860 7104 12872
rect 7156 12860 7162 12912
rect 6273 12835 6331 12841
rect 6273 12801 6285 12835
rect 6319 12801 6331 12835
rect 6273 12795 6331 12801
rect 8110 12792 8116 12844
rect 8168 12832 8174 12844
rect 8312 12832 8340 12940
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11885 12971 11943 12977
rect 11885 12937 11897 12971
rect 11931 12968 11943 12971
rect 12066 12968 12072 12980
rect 11931 12940 12072 12968
rect 11931 12937 11943 12940
rect 11885 12931 11943 12937
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 15286 12928 15292 12980
rect 15344 12928 15350 12980
rect 18141 12971 18199 12977
rect 18141 12937 18153 12971
rect 18187 12968 18199 12971
rect 18693 12971 18751 12977
rect 18693 12968 18705 12971
rect 18187 12940 18705 12968
rect 18187 12937 18199 12940
rect 18141 12931 18199 12937
rect 18693 12937 18705 12940
rect 18739 12937 18751 12971
rect 18693 12931 18751 12937
rect 20530 12928 20536 12980
rect 20588 12968 20594 12980
rect 20990 12968 20996 12980
rect 20588 12940 20996 12968
rect 20588 12928 20594 12940
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 21082 12928 21088 12980
rect 21140 12928 21146 12980
rect 21266 12928 21272 12980
rect 21324 12928 21330 12980
rect 21913 12971 21971 12977
rect 21913 12937 21925 12971
rect 21959 12968 21971 12971
rect 22741 12971 22799 12977
rect 22741 12968 22753 12971
rect 21959 12940 22753 12968
rect 21959 12937 21971 12940
rect 21913 12931 21971 12937
rect 22741 12937 22753 12940
rect 22787 12937 22799 12971
rect 22741 12931 22799 12937
rect 14918 12860 14924 12912
rect 14976 12900 14982 12912
rect 18509 12903 18567 12909
rect 14976 12872 16068 12900
rect 14976 12860 14982 12872
rect 8168 12804 8340 12832
rect 8168 12792 8174 12804
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10321 12835 10379 12841
rect 10321 12832 10333 12835
rect 10192 12804 10333 12832
rect 10192 12792 10198 12804
rect 10321 12801 10333 12804
rect 10367 12801 10379 12835
rect 10321 12795 10379 12801
rect 10520 12804 11744 12832
rect 5994 12724 6000 12776
rect 6052 12773 6058 12776
rect 6052 12764 6064 12773
rect 6365 12767 6423 12773
rect 6052 12736 6097 12764
rect 6052 12727 6064 12736
rect 6365 12733 6377 12767
rect 6411 12733 6423 12767
rect 6365 12727 6423 12733
rect 6052 12724 6058 12727
rect 6178 12656 6184 12708
rect 6236 12696 6242 12708
rect 6380 12696 6408 12727
rect 6546 12724 6552 12776
rect 6604 12724 6610 12776
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12764 7895 12767
rect 8386 12764 8392 12776
rect 7883 12736 8392 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12764 8631 12767
rect 8662 12764 8668 12776
rect 8619 12736 8668 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 10410 12724 10416 12776
rect 10468 12724 10474 12776
rect 6236 12668 6408 12696
rect 7929 12699 7987 12705
rect 6236 12656 6242 12668
rect 7929 12665 7941 12699
rect 7975 12696 7987 12699
rect 8478 12696 8484 12708
rect 7975 12668 8484 12696
rect 7975 12665 7987 12668
rect 7929 12659 7987 12665
rect 8478 12656 8484 12668
rect 8536 12656 8542 12708
rect 8840 12699 8898 12705
rect 8840 12665 8852 12699
rect 8886 12696 8898 12699
rect 9030 12696 9036 12708
rect 8886 12668 9036 12696
rect 8886 12665 8898 12668
rect 8840 12659 8898 12665
rect 9030 12656 9036 12668
rect 9088 12656 9094 12708
rect 9214 12656 9220 12708
rect 9272 12696 9278 12708
rect 10520 12696 10548 12804
rect 11716 12773 11744 12804
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 16040 12841 16068 12872
rect 18509 12869 18521 12903
rect 18555 12900 18567 12903
rect 19334 12900 19340 12912
rect 18555 12872 19340 12900
rect 18555 12869 18567 12872
rect 18509 12863 18567 12869
rect 19334 12860 19340 12872
rect 19392 12860 19398 12912
rect 22186 12860 22192 12912
rect 22244 12900 22250 12912
rect 22833 12903 22891 12909
rect 22833 12900 22845 12903
rect 22244 12872 22845 12900
rect 22244 12860 22250 12872
rect 22833 12869 22845 12872
rect 22879 12869 22891 12903
rect 22833 12863 22891 12869
rect 15841 12835 15899 12841
rect 15841 12832 15853 12835
rect 15620 12804 15853 12832
rect 15620 12792 15626 12804
rect 15841 12801 15853 12804
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12832 16083 12835
rect 16850 12832 16856 12844
rect 16071 12804 16856 12832
rect 16071 12801 16083 12804
rect 16025 12795 16083 12801
rect 16850 12792 16856 12804
rect 16908 12792 16914 12844
rect 18138 12832 18144 12844
rect 17696 12804 18144 12832
rect 11609 12767 11667 12773
rect 11609 12733 11621 12767
rect 11655 12733 11667 12767
rect 11609 12727 11667 12733
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12764 11759 12767
rect 12342 12764 12348 12776
rect 11747 12736 12348 12764
rect 11747 12733 11759 12736
rect 11701 12727 11759 12733
rect 9272 12668 10548 12696
rect 11624 12696 11652 12727
rect 12342 12724 12348 12736
rect 12400 12724 12406 12776
rect 12710 12724 12716 12776
rect 12768 12764 12774 12776
rect 13090 12767 13148 12773
rect 13090 12764 13102 12767
rect 12768 12736 13102 12764
rect 12768 12724 12774 12736
rect 13090 12733 13102 12736
rect 13136 12733 13148 12767
rect 13090 12727 13148 12733
rect 13354 12724 13360 12776
rect 13412 12724 13418 12776
rect 14182 12773 14188 12776
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12733 13967 12767
rect 14176 12764 14188 12773
rect 14143 12736 14188 12764
rect 13909 12727 13967 12733
rect 14176 12727 14188 12736
rect 12618 12696 12624 12708
rect 11624 12668 12624 12696
rect 9272 12656 9278 12668
rect 12618 12656 12624 12668
rect 12676 12656 12682 12708
rect 13924 12696 13952 12727
rect 14182 12724 14188 12727
rect 14240 12724 14246 12776
rect 17696 12773 17724 12804
rect 18138 12792 18144 12804
rect 18196 12832 18202 12844
rect 18196 12804 19196 12832
rect 18196 12792 18202 12804
rect 17681 12767 17739 12773
rect 17681 12733 17693 12767
rect 17727 12733 17739 12767
rect 17681 12727 17739 12733
rect 17862 12724 17868 12776
rect 17920 12764 17926 12776
rect 17920 12736 18552 12764
rect 17920 12724 17926 12736
rect 15470 12696 15476 12708
rect 13924 12668 15476 12696
rect 15470 12656 15476 12668
rect 15528 12656 15534 12708
rect 17773 12699 17831 12705
rect 17773 12665 17785 12699
rect 17819 12696 17831 12699
rect 18046 12696 18052 12708
rect 17819 12668 18052 12696
rect 17819 12665 17831 12668
rect 17773 12659 17831 12665
rect 18046 12656 18052 12668
rect 18104 12656 18110 12708
rect 18524 12696 18552 12736
rect 18598 12724 18604 12776
rect 18656 12764 18662 12776
rect 19168 12773 19196 12804
rect 18877 12767 18935 12773
rect 18877 12764 18889 12767
rect 18656 12736 18889 12764
rect 18656 12724 18662 12736
rect 18877 12733 18889 12736
rect 18923 12733 18935 12767
rect 18877 12727 18935 12733
rect 19153 12767 19211 12773
rect 19153 12733 19165 12767
rect 19199 12733 19211 12767
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19153 12727 19211 12733
rect 19352 12736 19625 12764
rect 19058 12696 19064 12708
rect 18524 12668 19064 12696
rect 19058 12656 19064 12668
rect 19116 12656 19122 12708
rect 19242 12656 19248 12708
rect 19300 12656 19306 12708
rect 4893 12631 4951 12637
rect 4893 12597 4905 12631
rect 4939 12628 4951 12631
rect 5534 12628 5540 12640
rect 4939 12600 5540 12628
rect 4939 12597 4951 12600
rect 4893 12591 4951 12597
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 6733 12631 6791 12637
rect 6733 12597 6745 12631
rect 6779 12628 6791 12631
rect 7098 12628 7104 12640
rect 6779 12600 7104 12628
rect 6779 12597 6791 12600
rect 6733 12591 6791 12597
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 9398 12628 9404 12640
rect 8996 12600 9404 12628
rect 8996 12588 9002 12600
rect 9398 12588 9404 12600
rect 9456 12628 9462 12640
rect 9953 12631 10011 12637
rect 9953 12628 9965 12631
rect 9456 12600 9965 12628
rect 9456 12588 9462 12600
rect 9953 12597 9965 12600
rect 9999 12597 10011 12631
rect 9953 12591 10011 12597
rect 10781 12631 10839 12637
rect 10781 12597 10793 12631
rect 10827 12628 10839 12631
rect 11698 12628 11704 12640
rect 10827 12600 11704 12628
rect 10827 12597 10839 12600
rect 10781 12591 10839 12597
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 11977 12631 12035 12637
rect 11977 12597 11989 12631
rect 12023 12628 12035 12631
rect 12526 12628 12532 12640
rect 12023 12600 12532 12628
rect 12023 12597 12035 12600
rect 11977 12591 12035 12597
rect 12526 12588 12532 12600
rect 12584 12628 12590 12640
rect 12710 12628 12716 12640
rect 12584 12600 12716 12628
rect 12584 12588 12590 12600
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 15378 12588 15384 12640
rect 15436 12588 15442 12640
rect 15746 12588 15752 12640
rect 15804 12588 15810 12640
rect 17954 12588 17960 12640
rect 18012 12588 18018 12640
rect 18141 12631 18199 12637
rect 18141 12597 18153 12631
rect 18187 12628 18199 12631
rect 18414 12628 18420 12640
rect 18187 12600 18420 12628
rect 18187 12597 18199 12600
rect 18141 12591 18199 12597
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 19150 12588 19156 12640
rect 19208 12628 19214 12640
rect 19352 12628 19380 12736
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 19702 12724 19708 12776
rect 19760 12764 19766 12776
rect 19869 12767 19927 12773
rect 19869 12764 19881 12767
rect 19760 12736 19881 12764
rect 19760 12724 19766 12736
rect 19869 12733 19881 12736
rect 19915 12733 19927 12767
rect 19869 12727 19927 12733
rect 21358 12724 21364 12776
rect 21416 12764 21422 12776
rect 21634 12764 21640 12776
rect 21416 12736 21640 12764
rect 21416 12724 21422 12736
rect 21634 12724 21640 12736
rect 21692 12764 21698 12776
rect 21692 12736 22094 12764
rect 21692 12724 21698 12736
rect 19426 12656 19432 12708
rect 19484 12696 19490 12708
rect 21269 12699 21327 12705
rect 21269 12696 21281 12699
rect 19484 12668 21281 12696
rect 19484 12656 19490 12668
rect 21269 12665 21281 12668
rect 21315 12696 21327 12699
rect 21450 12696 21456 12708
rect 21315 12668 21456 12696
rect 21315 12665 21327 12668
rect 21269 12659 21327 12665
rect 21450 12656 21456 12668
rect 21508 12656 21514 12708
rect 22066 12696 22094 12736
rect 22278 12724 22284 12776
rect 22336 12724 22342 12776
rect 23014 12724 23020 12776
rect 23072 12724 23078 12776
rect 22373 12699 22431 12705
rect 22373 12696 22385 12699
rect 22066 12668 22385 12696
rect 22373 12665 22385 12668
rect 22419 12665 22431 12699
rect 22373 12659 22431 12665
rect 22557 12699 22615 12705
rect 22557 12665 22569 12699
rect 22603 12696 22615 12699
rect 22922 12696 22928 12708
rect 22603 12668 22928 12696
rect 22603 12665 22615 12668
rect 22557 12659 22615 12665
rect 22922 12656 22928 12668
rect 22980 12656 22986 12708
rect 19208 12600 19380 12628
rect 19208 12588 19214 12600
rect 21726 12588 21732 12640
rect 21784 12588 21790 12640
rect 21910 12588 21916 12640
rect 21968 12588 21974 12640
rect 552 12538 23368 12560
rect 552 12486 4322 12538
rect 4374 12486 4386 12538
rect 4438 12486 4450 12538
rect 4502 12486 4514 12538
rect 4566 12486 4578 12538
rect 4630 12486 23368 12538
rect 552 12464 23368 12486
rect 5629 12427 5687 12433
rect 5629 12393 5641 12427
rect 5675 12424 5687 12427
rect 7190 12424 7196 12436
rect 5675 12396 7196 12424
rect 5675 12393 5687 12396
rect 5629 12387 5687 12393
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 11974 12424 11980 12436
rect 11204 12396 11980 12424
rect 11204 12384 11210 12396
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12618 12384 12624 12436
rect 12676 12424 12682 12436
rect 12713 12427 12771 12433
rect 12713 12424 12725 12427
rect 12676 12396 12725 12424
rect 12676 12384 12682 12396
rect 12713 12393 12725 12396
rect 12759 12393 12771 12427
rect 12713 12387 12771 12393
rect 13541 12427 13599 12433
rect 13541 12393 13553 12427
rect 13587 12424 13599 12427
rect 17862 12424 17868 12436
rect 13587 12396 14136 12424
rect 13587 12393 13599 12396
rect 13541 12387 13599 12393
rect 5534 12356 5540 12368
rect 5368 12328 5540 12356
rect 5368 12297 5396 12328
rect 5534 12316 5540 12328
rect 5592 12356 5598 12368
rect 5718 12356 5724 12368
rect 5592 12328 5724 12356
rect 5592 12316 5598 12328
rect 5718 12316 5724 12328
rect 5776 12356 5782 12368
rect 6457 12359 6515 12365
rect 5776 12328 6224 12356
rect 5776 12316 5782 12328
rect 6196 12297 6224 12328
rect 6457 12325 6469 12359
rect 6503 12356 6515 12359
rect 7006 12356 7012 12368
rect 6503 12328 7012 12356
rect 6503 12325 6515 12328
rect 6457 12319 6515 12325
rect 7006 12316 7012 12328
rect 7064 12356 7070 12368
rect 11606 12365 11612 12368
rect 11600 12356 11612 12365
rect 7064 12328 7328 12356
rect 11567 12328 11612 12356
rect 7064 12316 7070 12328
rect 5353 12291 5411 12297
rect 5353 12257 5365 12291
rect 5399 12257 5411 12291
rect 5353 12251 5411 12257
rect 5445 12291 5503 12297
rect 5445 12257 5457 12291
rect 5491 12288 5503 12291
rect 6181 12291 6239 12297
rect 5491 12260 6132 12288
rect 5491 12257 5503 12260
rect 5445 12251 5503 12257
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12189 5687 12223
rect 6104 12220 6132 12260
rect 6181 12257 6193 12291
rect 6227 12288 6239 12291
rect 6730 12288 6736 12300
rect 6227 12260 6736 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 7098 12248 7104 12300
rect 7156 12248 7162 12300
rect 7300 12297 7328 12328
rect 11600 12319 11612 12328
rect 11606 12316 11612 12319
rect 11664 12316 11670 12368
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12288 9275 12291
rect 10226 12288 10232 12300
rect 9263 12260 10232 12288
rect 9263 12257 9275 12260
rect 9217 12251 9275 12257
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 13354 12288 13360 12300
rect 11348 12260 13360 12288
rect 11348 12232 11376 12260
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12288 13783 12291
rect 13814 12288 13820 12300
rect 13771 12260 13820 12288
rect 13771 12257 13783 12260
rect 13725 12251 13783 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 13906 12248 13912 12300
rect 13964 12248 13970 12300
rect 14108 12288 14136 12396
rect 17420 12396 17868 12424
rect 16574 12316 16580 12368
rect 16632 12316 16638 12368
rect 17420 12365 17448 12396
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 18598 12384 18604 12436
rect 18656 12424 18662 12436
rect 19061 12427 19119 12433
rect 19061 12424 19073 12427
rect 18656 12396 19073 12424
rect 18656 12384 18662 12396
rect 19061 12393 19073 12396
rect 19107 12393 19119 12427
rect 19061 12387 19119 12393
rect 20625 12427 20683 12433
rect 20625 12393 20637 12427
rect 20671 12424 20683 12427
rect 20714 12424 20720 12436
rect 20671 12396 20720 12424
rect 20671 12393 20683 12396
rect 20625 12387 20683 12393
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 17954 12365 17960 12368
rect 17405 12359 17463 12365
rect 17405 12325 17417 12359
rect 17451 12325 17463 12359
rect 17948 12356 17960 12365
rect 17915 12328 17960 12356
rect 17405 12319 17463 12325
rect 17948 12319 17960 12328
rect 17954 12316 17960 12319
rect 18012 12316 18018 12368
rect 18138 12316 18144 12368
rect 18196 12316 18202 12368
rect 21726 12316 21732 12368
rect 21784 12356 21790 12368
rect 21882 12359 21940 12365
rect 21882 12356 21894 12359
rect 21784 12328 21894 12356
rect 21784 12316 21790 12328
rect 21882 12325 21894 12328
rect 21928 12325 21940 12359
rect 21882 12319 21940 12325
rect 14349 12291 14407 12297
rect 14349 12288 14361 12291
rect 14108 12260 14361 12288
rect 14349 12257 14361 12260
rect 14395 12257 14407 12291
rect 14349 12251 14407 12257
rect 16485 12291 16543 12297
rect 16485 12257 16497 12291
rect 16531 12288 16543 12291
rect 16592 12288 16620 12316
rect 16531 12260 16620 12288
rect 17589 12291 17647 12297
rect 16531 12257 16543 12260
rect 16485 12251 16543 12257
rect 17589 12257 17601 12291
rect 17635 12288 17647 12291
rect 18156 12288 18184 12316
rect 17635 12260 18184 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 18230 12248 18236 12300
rect 18288 12288 18294 12300
rect 19409 12291 19467 12297
rect 19409 12288 19421 12291
rect 18288 12260 19421 12288
rect 18288 12248 18294 12260
rect 19409 12257 19421 12260
rect 19455 12257 19467 12291
rect 19409 12251 19467 12257
rect 20806 12248 20812 12300
rect 20864 12248 20870 12300
rect 20990 12248 20996 12300
rect 21048 12248 21054 12300
rect 21082 12248 21088 12300
rect 21140 12288 21146 12300
rect 21361 12291 21419 12297
rect 21361 12288 21373 12291
rect 21140 12260 21373 12288
rect 21140 12248 21146 12260
rect 21361 12257 21373 12260
rect 21407 12288 21419 12291
rect 22646 12288 22652 12300
rect 21407 12260 22652 12288
rect 21407 12257 21419 12260
rect 21361 12251 21419 12257
rect 22646 12248 22652 12260
rect 22704 12248 22710 12300
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 6104 12192 6285 12220
rect 5629 12183 5687 12189
rect 6273 12189 6285 12192
rect 6319 12220 6331 12223
rect 6362 12220 6368 12232
rect 6319 12192 6368 12220
rect 6319 12189 6331 12192
rect 6273 12183 6331 12189
rect 5644 12152 5672 12183
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 6178 12152 6184 12164
rect 5644 12124 6184 12152
rect 6178 12112 6184 12124
rect 6236 12152 6242 12164
rect 6564 12152 6592 12183
rect 9306 12180 9312 12232
rect 9364 12180 9370 12232
rect 11330 12180 11336 12232
rect 11388 12180 11394 12232
rect 14001 12223 14059 12229
rect 14001 12189 14013 12223
rect 14047 12189 14059 12223
rect 14001 12183 14059 12189
rect 6236 12124 6592 12152
rect 6917 12155 6975 12161
rect 6236 12112 6242 12124
rect 6917 12121 6929 12155
rect 6963 12152 6975 12155
rect 7466 12152 7472 12164
rect 6963 12124 7472 12152
rect 6963 12121 6975 12124
rect 6917 12115 6975 12121
rect 7466 12112 7472 12124
rect 7524 12112 7530 12164
rect 5810 12044 5816 12096
rect 5868 12044 5874 12096
rect 6362 12044 6368 12096
rect 6420 12084 6426 12096
rect 6457 12087 6515 12093
rect 6457 12084 6469 12087
rect 6420 12056 6469 12084
rect 6420 12044 6426 12056
rect 6457 12053 6469 12056
rect 6503 12053 6515 12087
rect 6457 12047 6515 12053
rect 7193 12087 7251 12093
rect 7193 12053 7205 12087
rect 7239 12084 7251 12087
rect 7374 12084 7380 12096
rect 7239 12056 7380 12084
rect 7239 12053 7251 12056
rect 7193 12047 7251 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 9493 12087 9551 12093
rect 9493 12053 9505 12087
rect 9539 12084 9551 12087
rect 9858 12084 9864 12096
rect 9539 12056 9864 12084
rect 9539 12053 9551 12056
rect 9493 12047 9551 12053
rect 9858 12044 9864 12056
rect 9916 12044 9922 12096
rect 14016 12084 14044 12183
rect 14090 12180 14096 12232
rect 14148 12180 14154 12232
rect 16574 12180 16580 12232
rect 16632 12220 16638 12232
rect 16758 12220 16764 12232
rect 16632 12192 16764 12220
rect 16632 12180 16638 12192
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12189 17739 12223
rect 17681 12183 17739 12189
rect 15102 12112 15108 12164
rect 15160 12152 15166 12164
rect 17696 12152 17724 12183
rect 19150 12180 19156 12232
rect 19208 12180 19214 12232
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 21637 12223 21695 12229
rect 21637 12220 21649 12223
rect 21324 12192 21649 12220
rect 21324 12180 21330 12192
rect 21637 12189 21649 12192
rect 21683 12189 21695 12223
rect 21637 12183 21695 12189
rect 15160 12124 17724 12152
rect 15160 12112 15166 12124
rect 14826 12084 14832 12096
rect 14016 12056 14832 12084
rect 14826 12044 14832 12056
rect 14884 12084 14890 12096
rect 15473 12087 15531 12093
rect 15473 12084 15485 12087
rect 14884 12056 15485 12084
rect 14884 12044 14890 12056
rect 15473 12053 15485 12056
rect 15519 12084 15531 12087
rect 16114 12084 16120 12096
rect 15519 12056 16120 12084
rect 15519 12053 15531 12056
rect 15473 12047 15531 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16850 12044 16856 12096
rect 16908 12044 16914 12096
rect 17221 12087 17279 12093
rect 17221 12053 17233 12087
rect 17267 12084 17279 12087
rect 17954 12084 17960 12096
rect 17267 12056 17960 12084
rect 17267 12053 17279 12056
rect 17221 12047 17279 12053
rect 17954 12044 17960 12056
rect 18012 12044 18018 12096
rect 19058 12044 19064 12096
rect 19116 12084 19122 12096
rect 20533 12087 20591 12093
rect 20533 12084 20545 12087
rect 19116 12056 20545 12084
rect 19116 12044 19122 12056
rect 20533 12053 20545 12056
rect 20579 12053 20591 12087
rect 20533 12047 20591 12053
rect 21450 12044 21456 12096
rect 21508 12084 21514 12096
rect 21634 12084 21640 12096
rect 21508 12056 21640 12084
rect 21508 12044 21514 12056
rect 21634 12044 21640 12056
rect 21692 12084 21698 12096
rect 21910 12084 21916 12096
rect 21692 12056 21916 12084
rect 21692 12044 21698 12056
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 22922 12044 22928 12096
rect 22980 12084 22986 12096
rect 23017 12087 23075 12093
rect 23017 12084 23029 12087
rect 22980 12056 23029 12084
rect 22980 12044 22986 12056
rect 23017 12053 23029 12056
rect 23063 12053 23075 12087
rect 23017 12047 23075 12053
rect 552 11994 23368 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 23368 11994
rect 552 11920 23368 11942
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 7098 11880 7104 11892
rect 6687 11852 7104 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 16025 11883 16083 11889
rect 16025 11880 16037 11883
rect 15804 11852 16037 11880
rect 15804 11840 15810 11852
rect 16025 11849 16037 11852
rect 16071 11849 16083 11883
rect 16025 11843 16083 11849
rect 6914 11772 6920 11824
rect 6972 11772 6978 11824
rect 5810 11704 5816 11756
rect 5868 11744 5874 11756
rect 5905 11747 5963 11753
rect 5905 11744 5917 11747
rect 5868 11716 5917 11744
rect 5868 11704 5874 11716
rect 5905 11713 5917 11716
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 6696 11716 7236 11744
rect 6696 11704 6702 11716
rect 7208 11688 7236 11716
rect 7466 11704 7472 11756
rect 7524 11744 7530 11756
rect 8294 11744 8300 11756
rect 7524 11716 8300 11744
rect 7524 11704 7530 11716
rect 8294 11704 8300 11716
rect 8352 11744 8358 11756
rect 8573 11747 8631 11753
rect 8573 11744 8585 11747
rect 8352 11716 8585 11744
rect 8352 11704 8358 11716
rect 8573 11713 8585 11716
rect 8619 11713 8631 11747
rect 8573 11707 8631 11713
rect 5994 11636 6000 11688
rect 6052 11636 6058 11688
rect 6472 11648 6868 11676
rect 6472 11620 6500 11648
rect 6454 11568 6460 11620
rect 6512 11568 6518 11620
rect 6840 11608 6868 11648
rect 7098 11636 7104 11688
rect 7156 11636 7162 11688
rect 7190 11636 7196 11688
rect 7248 11636 7254 11688
rect 8386 11636 8392 11688
rect 8444 11676 8450 11688
rect 8481 11679 8539 11685
rect 8481 11676 8493 11679
rect 8444 11648 8493 11676
rect 8444 11636 8450 11648
rect 8481 11645 8493 11648
rect 8527 11645 8539 11679
rect 8481 11639 8539 11645
rect 6917 11611 6975 11617
rect 6917 11608 6929 11611
rect 6840 11580 6929 11608
rect 6917 11577 6929 11580
rect 6963 11577 6975 11611
rect 8588 11608 8616 11707
rect 8754 11704 8760 11756
rect 8812 11704 8818 11756
rect 16040 11744 16068 11843
rect 16114 11840 16120 11892
rect 16172 11840 16178 11892
rect 16574 11840 16580 11892
rect 16632 11840 16638 11892
rect 16758 11840 16764 11892
rect 16816 11880 16822 11892
rect 17037 11883 17095 11889
rect 17037 11880 17049 11883
rect 16816 11852 17049 11880
rect 16816 11840 16822 11852
rect 17037 11849 17049 11852
rect 17083 11849 17095 11883
rect 17037 11843 17095 11849
rect 18046 11840 18052 11892
rect 18104 11840 18110 11892
rect 18230 11840 18236 11892
rect 18288 11840 18294 11892
rect 19429 11883 19487 11889
rect 19429 11849 19441 11883
rect 19475 11880 19487 11883
rect 20346 11880 20352 11892
rect 19475 11852 20352 11880
rect 19475 11849 19487 11852
rect 19429 11843 19487 11849
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 21085 11883 21143 11889
rect 21085 11849 21097 11883
rect 21131 11880 21143 11883
rect 21174 11880 21180 11892
rect 21131 11852 21180 11880
rect 21131 11849 21143 11852
rect 21085 11843 21143 11849
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 21545 11883 21603 11889
rect 21545 11849 21557 11883
rect 21591 11880 21603 11883
rect 22278 11880 22284 11892
rect 21591 11852 22284 11880
rect 21591 11849 21603 11852
rect 21545 11843 21603 11849
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 17497 11815 17555 11821
rect 17497 11781 17509 11815
rect 17543 11812 17555 11815
rect 18782 11812 18788 11824
rect 17543 11784 18788 11812
rect 17543 11781 17555 11784
rect 17497 11775 17555 11781
rect 18782 11772 18788 11784
rect 18840 11772 18846 11824
rect 16209 11747 16267 11753
rect 16209 11744 16221 11747
rect 16040 11716 16221 11744
rect 16209 11713 16221 11716
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 21177 11747 21235 11753
rect 21177 11713 21189 11747
rect 21223 11744 21235 11747
rect 21223 11716 21772 11744
rect 21223 11713 21235 11716
rect 21177 11707 21235 11713
rect 8662 11636 8668 11688
rect 8720 11676 8726 11688
rect 8849 11679 8907 11685
rect 8849 11676 8861 11679
rect 8720 11648 8861 11676
rect 8720 11636 8726 11648
rect 8849 11645 8861 11648
rect 8895 11645 8907 11679
rect 10226 11676 10232 11688
rect 8849 11639 8907 11645
rect 9048 11648 10232 11676
rect 9048 11608 9076 11648
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 10965 11679 11023 11685
rect 10965 11645 10977 11679
rect 11011 11676 11023 11679
rect 11011 11648 11376 11676
rect 11011 11645 11023 11648
rect 10965 11639 11023 11645
rect 11348 11620 11376 11648
rect 14090 11636 14096 11688
rect 14148 11676 14154 11688
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 14148 11648 14657 11676
rect 14148 11636 14154 11648
rect 14645 11645 14657 11648
rect 14691 11645 14703 11679
rect 14645 11639 14703 11645
rect 14912 11679 14970 11685
rect 14912 11645 14924 11679
rect 14958 11676 14970 11679
rect 15378 11676 15384 11688
rect 14958 11648 15384 11676
rect 14958 11645 14970 11648
rect 14912 11639 14970 11645
rect 8588 11580 9076 11608
rect 9116 11611 9174 11617
rect 6917 11571 6975 11577
rect 9116 11577 9128 11611
rect 9162 11608 9174 11611
rect 9398 11608 9404 11620
rect 9162 11580 9404 11608
rect 9162 11577 9174 11580
rect 9116 11571 9174 11577
rect 9398 11568 9404 11580
rect 9456 11568 9462 11620
rect 11238 11617 11244 11620
rect 11232 11571 11244 11617
rect 11238 11568 11244 11571
rect 11296 11568 11302 11620
rect 11330 11568 11336 11620
rect 11388 11568 11394 11620
rect 14660 11608 14688 11639
rect 15378 11636 15384 11648
rect 15436 11636 15442 11688
rect 16393 11679 16451 11685
rect 16393 11676 16405 11679
rect 15488 11648 16405 11676
rect 15010 11608 15016 11620
rect 14660 11580 15016 11608
rect 15010 11568 15016 11580
rect 15068 11568 15074 11620
rect 15194 11568 15200 11620
rect 15252 11608 15258 11620
rect 15488 11608 15516 11648
rect 16393 11645 16405 11648
rect 16439 11645 16451 11679
rect 16393 11639 16451 11645
rect 17218 11636 17224 11688
rect 17276 11636 17282 11688
rect 17313 11679 17371 11685
rect 17313 11645 17325 11679
rect 17359 11676 17371 11679
rect 17402 11676 17408 11688
rect 17359 11648 17408 11676
rect 17359 11645 17371 11648
rect 17313 11639 17371 11645
rect 17402 11636 17408 11648
rect 17460 11636 17466 11688
rect 19426 11676 19432 11688
rect 17880 11648 19432 11676
rect 15252 11580 15516 11608
rect 16117 11611 16175 11617
rect 15252 11568 15258 11580
rect 16117 11577 16129 11611
rect 16163 11577 16175 11611
rect 16117 11571 16175 11577
rect 6365 11543 6423 11549
rect 6365 11509 6377 11543
rect 6411 11540 6423 11543
rect 6546 11540 6552 11552
rect 6411 11512 6552 11540
rect 6411 11509 6423 11512
rect 6365 11503 6423 11509
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 6638 11500 6644 11552
rect 6696 11549 6702 11552
rect 6696 11543 6715 11549
rect 6703 11509 6715 11543
rect 6696 11503 6715 11509
rect 6696 11500 6702 11503
rect 6822 11500 6828 11552
rect 6880 11500 6886 11552
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 8570 11540 8576 11552
rect 7708 11512 8576 11540
rect 7708 11500 7714 11512
rect 8570 11500 8576 11512
rect 8628 11500 8634 11552
rect 8757 11543 8815 11549
rect 8757 11509 8769 11543
rect 8803 11540 8815 11543
rect 9214 11540 9220 11552
rect 8803 11512 9220 11540
rect 8803 11509 8815 11512
rect 8757 11503 8815 11509
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 10229 11543 10287 11549
rect 10229 11509 10241 11543
rect 10275 11540 10287 11543
rect 10318 11540 10324 11552
rect 10275 11512 10324 11540
rect 10275 11509 10287 11512
rect 10229 11503 10287 11509
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 12342 11500 12348 11552
rect 12400 11500 12406 11552
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 16132 11540 16160 11571
rect 16666 11568 16672 11620
rect 16724 11608 16730 11620
rect 17880 11617 17908 11648
rect 19426 11636 19432 11648
rect 19484 11636 19490 11688
rect 19705 11679 19763 11685
rect 19705 11645 19717 11679
rect 19751 11676 19763 11679
rect 19751 11648 21312 11676
rect 19751 11645 19763 11648
rect 19705 11639 19763 11645
rect 21284 11620 21312 11648
rect 21358 11636 21364 11688
rect 21416 11636 21422 11688
rect 21637 11679 21695 11685
rect 21637 11676 21649 11679
rect 21468 11648 21649 11676
rect 17037 11611 17095 11617
rect 17037 11608 17049 11611
rect 16724 11580 17049 11608
rect 16724 11568 16730 11580
rect 17037 11577 17049 11580
rect 17083 11577 17095 11611
rect 17037 11571 17095 11577
rect 17865 11611 17923 11617
rect 17865 11577 17877 11611
rect 17911 11577 17923 11611
rect 17865 11571 17923 11577
rect 15344 11512 16160 11540
rect 15344 11500 15350 11512
rect 17310 11500 17316 11552
rect 17368 11540 17374 11552
rect 17880 11540 17908 11571
rect 17954 11568 17960 11620
rect 18012 11608 18018 11620
rect 18065 11611 18123 11617
rect 18065 11608 18077 11611
rect 18012 11580 18077 11608
rect 18012 11568 18018 11580
rect 18065 11577 18077 11580
rect 18111 11577 18123 11611
rect 18065 11571 18123 11577
rect 18414 11568 18420 11620
rect 18472 11608 18478 11620
rect 19245 11611 19303 11617
rect 19245 11608 19257 11611
rect 18472 11580 19257 11608
rect 18472 11568 18478 11580
rect 19245 11577 19257 11580
rect 19291 11608 19303 11611
rect 19334 11608 19340 11620
rect 19291 11580 19340 11608
rect 19291 11577 19303 11580
rect 19245 11571 19303 11577
rect 19334 11568 19340 11580
rect 19392 11568 19398 11620
rect 19950 11611 20008 11617
rect 19950 11608 19962 11611
rect 19628 11580 19962 11608
rect 17368 11512 17908 11540
rect 17368 11500 17374 11512
rect 19426 11500 19432 11552
rect 19484 11549 19490 11552
rect 19628 11549 19656 11580
rect 19950 11577 19962 11580
rect 19996 11577 20008 11611
rect 19950 11571 20008 11577
rect 21266 11568 21272 11620
rect 21324 11608 21330 11620
rect 21468 11608 21496 11648
rect 21637 11645 21649 11648
rect 21683 11645 21695 11679
rect 21744 11676 21772 11716
rect 22922 11676 22928 11688
rect 21744 11648 22928 11676
rect 21637 11639 21695 11645
rect 22922 11636 22928 11648
rect 22980 11636 22986 11688
rect 21324 11580 21496 11608
rect 21324 11568 21330 11580
rect 21542 11568 21548 11620
rect 21600 11608 21606 11620
rect 21882 11611 21940 11617
rect 21882 11608 21894 11611
rect 21600 11580 21894 11608
rect 21600 11568 21606 11580
rect 21882 11577 21894 11580
rect 21928 11577 21940 11611
rect 21882 11571 21940 11577
rect 19484 11543 19503 11549
rect 19491 11509 19503 11543
rect 19484 11503 19503 11509
rect 19613 11543 19671 11549
rect 19613 11509 19625 11543
rect 19659 11509 19671 11543
rect 19613 11503 19671 11509
rect 19484 11500 19490 11503
rect 22370 11500 22376 11552
rect 22428 11540 22434 11552
rect 23017 11543 23075 11549
rect 23017 11540 23029 11543
rect 22428 11512 23029 11540
rect 22428 11500 22434 11512
rect 23017 11509 23029 11512
rect 23063 11509 23075 11543
rect 23017 11503 23075 11509
rect 552 11450 23368 11472
rect 552 11398 4322 11450
rect 4374 11398 4386 11450
rect 4438 11398 4450 11450
rect 4502 11398 4514 11450
rect 4566 11398 4578 11450
rect 4630 11398 23368 11450
rect 552 11376 23368 11398
rect 5471 11339 5529 11345
rect 5471 11305 5483 11339
rect 5517 11336 5529 11339
rect 7101 11339 7159 11345
rect 7101 11336 7113 11339
rect 5517 11308 7113 11336
rect 5517 11305 5529 11308
rect 5471 11299 5529 11305
rect 7101 11305 7113 11308
rect 7147 11305 7159 11339
rect 7101 11299 7159 11305
rect 7466 11296 7472 11348
rect 7524 11296 7530 11348
rect 8113 11339 8171 11345
rect 8113 11305 8125 11339
rect 8159 11336 8171 11339
rect 9306 11336 9312 11348
rect 8159 11308 9312 11336
rect 8159 11305 8171 11308
rect 8113 11299 8171 11305
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 9398 11296 9404 11348
rect 9456 11296 9462 11348
rect 9858 11296 9864 11348
rect 9916 11296 9922 11348
rect 10689 11339 10747 11345
rect 10689 11305 10701 11339
rect 10735 11305 10747 11339
rect 10689 11299 10747 11305
rect 5261 11271 5319 11277
rect 5261 11237 5273 11271
rect 5307 11268 5319 11271
rect 5626 11268 5632 11280
rect 5307 11240 5632 11268
rect 5307 11237 5319 11240
rect 5261 11231 5319 11237
rect 5626 11228 5632 11240
rect 5684 11268 5690 11280
rect 5684 11240 6132 11268
rect 5684 11228 5690 11240
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11200 5227 11203
rect 5718 11200 5724 11212
rect 5215 11172 5724 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 4614 11092 4620 11144
rect 4672 11132 4678 11144
rect 5000 11132 5028 11163
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 5810 11160 5816 11212
rect 5868 11160 5874 11212
rect 5994 11160 6000 11212
rect 6052 11160 6058 11212
rect 6104 11200 6132 11240
rect 6178 11228 6184 11280
rect 6236 11228 6242 11280
rect 6365 11271 6423 11277
rect 6365 11237 6377 11271
rect 6411 11268 6423 11271
rect 6411 11240 6500 11268
rect 6411 11237 6423 11240
rect 6365 11231 6423 11237
rect 6273 11203 6331 11209
rect 6273 11200 6285 11203
rect 6104 11172 6285 11200
rect 6273 11169 6285 11172
rect 6319 11169 6331 11203
rect 6273 11163 6331 11169
rect 5074 11132 5080 11144
rect 4672 11104 5080 11132
rect 4672 11092 4678 11104
rect 5074 11092 5080 11104
rect 5132 11132 5138 11144
rect 6178 11132 6184 11144
rect 5132 11104 6184 11132
rect 5132 11092 5138 11104
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 4801 10999 4859 11005
rect 4801 10965 4813 10999
rect 4847 10996 4859 10999
rect 5445 10999 5503 11005
rect 5445 10996 5457 10999
rect 4847 10968 5457 10996
rect 4847 10965 4859 10968
rect 4801 10959 4859 10965
rect 5445 10965 5457 10968
rect 5491 10965 5503 10999
rect 5445 10959 5503 10965
rect 5629 10999 5687 11005
rect 5629 10965 5641 10999
rect 5675 10996 5687 10999
rect 6472 10996 6500 11240
rect 6730 11228 6736 11280
rect 6788 11268 6794 11280
rect 8357 11271 8415 11277
rect 8357 11268 8369 11271
rect 6788 11240 7328 11268
rect 6788 11228 6794 11240
rect 6546 11160 6552 11212
rect 6604 11200 6610 11212
rect 6641 11203 6699 11209
rect 6641 11200 6653 11203
rect 6604 11172 6653 11200
rect 6604 11160 6610 11172
rect 6641 11169 6653 11172
rect 6687 11169 6699 11203
rect 6641 11163 6699 11169
rect 6822 11160 6828 11212
rect 6880 11160 6886 11212
rect 7098 11160 7104 11212
rect 7156 11160 7162 11212
rect 7300 11209 7328 11240
rect 7392 11240 8369 11268
rect 7392 11212 7420 11240
rect 8357 11237 8369 11240
rect 8403 11237 8415 11271
rect 8357 11231 8415 11237
rect 8570 11228 8576 11280
rect 8628 11228 8634 11280
rect 9048 11240 10548 11268
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7374 11160 7380 11212
rect 7432 11160 7438 11212
rect 7650 11160 7656 11212
rect 7708 11160 7714 11212
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11169 7803 11203
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 7745 11163 7803 11169
rect 8312 11172 8953 11200
rect 7760 11132 7788 11163
rect 8312 11144 8340 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 7024 11104 7788 11132
rect 7837 11135 7895 11141
rect 7024 11073 7052 11104
rect 7837 11101 7849 11135
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 7009 11067 7067 11073
rect 7009 11033 7021 11067
rect 7055 11033 7067 11067
rect 7852 11064 7880 11095
rect 8294 11092 8300 11144
rect 8352 11092 8358 11144
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 9048 11141 9076 11240
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11200 9827 11203
rect 9815 11172 10088 11200
rect 9815 11169 9827 11172
rect 9769 11163 9827 11169
rect 9033 11135 9091 11141
rect 9033 11132 9045 11135
rect 8444 11104 9045 11132
rect 8444 11092 8450 11104
rect 9033 11101 9045 11104
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11101 10011 11135
rect 10060 11132 10088 11172
rect 10226 11160 10232 11212
rect 10284 11160 10290 11212
rect 10520 11209 10548 11240
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11169 10563 11203
rect 10704 11200 10732 11299
rect 11238 11296 11244 11348
rect 11296 11296 11302 11348
rect 11698 11296 11704 11348
rect 11756 11296 11762 11348
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11336 15531 11339
rect 16593 11339 16651 11345
rect 16593 11336 16605 11339
rect 15519 11308 16605 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 10980 11240 12296 11268
rect 10980 11209 11008 11240
rect 12268 11209 12296 11240
rect 14292 11240 15332 11268
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 10704 11172 10977 11200
rect 10505 11163 10563 11169
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11200 11207 11203
rect 11609 11203 11667 11209
rect 11609 11200 11621 11203
rect 11195 11172 11621 11200
rect 11195 11169 11207 11172
rect 11149 11163 11207 11169
rect 11609 11169 11621 11172
rect 11655 11200 11667 11203
rect 12253 11203 12311 11209
rect 11655 11172 12020 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 10318 11132 10324 11144
rect 10060 11104 10324 11132
rect 9953 11095 10011 11101
rect 8205 11067 8263 11073
rect 8205 11064 8217 11067
rect 7852 11036 8217 11064
rect 7009 11027 7067 11033
rect 8205 11033 8217 11036
rect 8251 11033 8263 11067
rect 8205 11027 8263 11033
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 9968 11064 9996 11095
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 11054 11092 11060 11144
rect 11112 11092 11118 11144
rect 11793 11135 11851 11141
rect 11793 11132 11805 11135
rect 11256 11104 11805 11132
rect 8812 11036 9628 11064
rect 9968 11036 10364 11064
rect 8812 11024 8818 11036
rect 5675 10968 6500 10996
rect 6825 10999 6883 11005
rect 5675 10965 5687 10968
rect 5629 10959 5687 10965
rect 6825 10965 6837 10999
rect 6871 10996 6883 10999
rect 6914 10996 6920 11008
rect 6871 10968 6920 10996
rect 6871 10965 6883 10968
rect 6825 10959 6883 10965
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 7653 10999 7711 11005
rect 7653 10965 7665 10999
rect 7699 10996 7711 10999
rect 7745 10999 7803 11005
rect 7745 10996 7757 10999
rect 7699 10968 7757 10996
rect 7699 10965 7711 10968
rect 7653 10959 7711 10965
rect 7745 10965 7757 10968
rect 7791 10965 7803 10999
rect 7745 10959 7803 10965
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 9140 11005 9168 11036
rect 8389 10999 8447 11005
rect 8389 10996 8401 10999
rect 8352 10968 8401 10996
rect 8352 10956 8358 10968
rect 8389 10965 8401 10968
rect 8435 10965 8447 10999
rect 8389 10959 8447 10965
rect 9125 10999 9183 11005
rect 9125 10965 9137 10999
rect 9171 10965 9183 10999
rect 9125 10959 9183 10965
rect 9309 10999 9367 11005
rect 9309 10965 9321 10999
rect 9355 10996 9367 10999
rect 9490 10996 9496 11008
rect 9355 10968 9496 10996
rect 9355 10965 9367 10968
rect 9309 10959 9367 10965
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 9600 10996 9628 11036
rect 10229 10999 10287 11005
rect 10229 10996 10241 10999
rect 9600 10968 10241 10996
rect 10229 10965 10241 10968
rect 10275 10965 10287 10999
rect 10336 10996 10364 11036
rect 11146 10996 11152 11008
rect 10336 10968 11152 10996
rect 10229 10959 10287 10965
rect 11146 10956 11152 10968
rect 11204 10996 11210 11008
rect 11256 10996 11284 11104
rect 11793 11101 11805 11104
rect 11839 11101 11851 11135
rect 11992 11132 12020 11172
rect 12253 11169 12265 11203
rect 12299 11200 12311 11203
rect 12526 11200 12532 11212
rect 12299 11172 12532 11200
rect 12299 11169 12311 11172
rect 12253 11163 12311 11169
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 12710 11160 12716 11212
rect 12768 11160 12774 11212
rect 12805 11203 12863 11209
rect 12805 11169 12817 11203
rect 12851 11169 12863 11203
rect 12805 11163 12863 11169
rect 12342 11132 12348 11144
rect 11992 11104 12348 11132
rect 11793 11095 11851 11101
rect 12342 11092 12348 11104
rect 12400 11132 12406 11144
rect 12437 11135 12495 11141
rect 12437 11132 12449 11135
rect 12400 11104 12449 11132
rect 12400 11092 12406 11104
rect 12437 11101 12449 11104
rect 12483 11132 12495 11135
rect 12820 11132 12848 11163
rect 13722 11160 13728 11212
rect 13780 11200 13786 11212
rect 14292 11209 14320 11240
rect 14752 11209 14780 11240
rect 15304 11212 15332 11240
rect 14277 11203 14335 11209
rect 14277 11200 14289 11203
rect 13780 11172 14289 11200
rect 13780 11160 13786 11172
rect 14277 11169 14289 11172
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11200 14519 11203
rect 14737 11203 14795 11209
rect 14507 11172 14596 11200
rect 14507 11169 14519 11172
rect 14461 11163 14519 11169
rect 14568 11141 14596 11172
rect 14737 11169 14749 11203
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 15013 11203 15071 11209
rect 15013 11169 15025 11203
rect 15059 11200 15071 11203
rect 15194 11200 15200 11212
rect 15059 11172 15200 11200
rect 15059 11169 15071 11172
rect 15013 11163 15071 11169
rect 12483 11104 12848 11132
rect 14553 11135 14611 11141
rect 12483 11101 12495 11104
rect 12437 11095 12495 11101
rect 14553 11101 14565 11135
rect 14599 11132 14611 11135
rect 15028 11132 15056 11163
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 15286 11160 15292 11212
rect 15344 11160 15350 11212
rect 15473 11203 15531 11209
rect 15473 11169 15485 11203
rect 15519 11200 15531 11203
rect 15562 11200 15568 11212
rect 15519 11172 15568 11200
rect 15519 11169 15531 11172
rect 15473 11163 15531 11169
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 15672 11209 15700 11308
rect 16593 11305 16605 11308
rect 16639 11305 16651 11339
rect 16593 11299 16651 11305
rect 16758 11296 16764 11348
rect 16816 11296 16822 11348
rect 17402 11296 17408 11348
rect 17460 11296 17466 11348
rect 17586 11296 17592 11348
rect 17644 11336 17650 11348
rect 17773 11339 17831 11345
rect 17773 11336 17785 11339
rect 17644 11308 17785 11336
rect 17644 11296 17650 11308
rect 17773 11305 17785 11308
rect 17819 11305 17831 11339
rect 17773 11299 17831 11305
rect 18049 11339 18107 11345
rect 18049 11305 18061 11339
rect 18095 11336 18107 11339
rect 18138 11336 18144 11348
rect 18095 11308 18144 11336
rect 18095 11305 18107 11308
rect 18049 11299 18107 11305
rect 18138 11296 18144 11308
rect 18196 11336 18202 11348
rect 18196 11308 18736 11336
rect 18196 11296 18202 11308
rect 15933 11271 15991 11277
rect 15933 11237 15945 11271
rect 15979 11268 15991 11271
rect 16390 11268 16396 11280
rect 15979 11240 16396 11268
rect 15979 11237 15991 11240
rect 15933 11231 15991 11237
rect 16390 11228 16396 11240
rect 16448 11268 16454 11280
rect 17497 11271 17555 11277
rect 17497 11268 17509 11271
rect 16448 11240 17509 11268
rect 16448 11228 16454 11240
rect 17497 11237 17509 11240
rect 17543 11237 17555 11271
rect 17497 11231 17555 11237
rect 18325 11271 18383 11277
rect 18325 11237 18337 11271
rect 18371 11268 18383 11271
rect 18414 11268 18420 11280
rect 18371 11240 18420 11268
rect 18371 11237 18383 11240
rect 18325 11231 18383 11237
rect 18414 11228 18420 11240
rect 18472 11228 18478 11280
rect 15657 11203 15715 11209
rect 15657 11169 15669 11203
rect 15703 11169 15715 11203
rect 15657 11163 15715 11169
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11169 15807 11203
rect 15749 11163 15807 11169
rect 14599 11104 15056 11132
rect 15764 11132 15792 11163
rect 17034 11160 17040 11212
rect 17092 11200 17098 11212
rect 17681 11203 17739 11209
rect 17681 11200 17693 11203
rect 17092 11172 17693 11200
rect 17092 11160 17098 11172
rect 17681 11169 17693 11172
rect 17727 11169 17739 11203
rect 17681 11163 17739 11169
rect 17862 11160 17868 11212
rect 17920 11160 17926 11212
rect 18708 11209 18736 11308
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 20073 11339 20131 11345
rect 20073 11336 20085 11339
rect 19484 11308 20085 11336
rect 19484 11296 19490 11308
rect 20073 11305 20085 11308
rect 20119 11305 20131 11339
rect 20073 11299 20131 11305
rect 20346 11296 20352 11348
rect 20404 11336 20410 11348
rect 20533 11339 20591 11345
rect 20533 11336 20545 11339
rect 20404 11308 20545 11336
rect 20404 11296 20410 11308
rect 20533 11305 20545 11308
rect 20579 11305 20591 11339
rect 20533 11299 20591 11305
rect 21542 11296 21548 11348
rect 21600 11296 21606 11348
rect 21634 11296 21640 11348
rect 21692 11336 21698 11348
rect 21729 11339 21787 11345
rect 21729 11336 21741 11339
rect 21692 11308 21741 11336
rect 21692 11296 21698 11308
rect 21729 11305 21741 11308
rect 21775 11305 21787 11339
rect 21729 11299 21787 11305
rect 20441 11271 20499 11277
rect 20441 11237 20453 11271
rect 20487 11268 20499 11271
rect 20487 11240 20760 11268
rect 20487 11237 20499 11240
rect 20441 11231 20499 11237
rect 20732 11212 20760 11240
rect 22278 11228 22284 11280
rect 22336 11268 22342 11280
rect 22557 11271 22615 11277
rect 22557 11268 22569 11271
rect 22336 11240 22569 11268
rect 22336 11228 22342 11240
rect 22557 11237 22569 11240
rect 22603 11237 22615 11271
rect 22557 11231 22615 11237
rect 18693 11203 18751 11209
rect 18693 11169 18705 11203
rect 18739 11169 18751 11203
rect 18693 11163 18751 11169
rect 20257 11203 20315 11209
rect 20257 11169 20269 11203
rect 20303 11200 20315 11203
rect 20533 11203 20591 11209
rect 20533 11200 20545 11203
rect 20303 11172 20545 11200
rect 20303 11169 20315 11172
rect 20257 11163 20315 11169
rect 20533 11169 20545 11172
rect 20579 11169 20591 11203
rect 20533 11163 20591 11169
rect 16574 11132 16580 11144
rect 15764 11104 16580 11132
rect 14599 11101 14611 11104
rect 14553 11095 14611 11101
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 16945 11135 17003 11141
rect 16945 11132 16957 11135
rect 16908 11104 16957 11132
rect 16908 11092 16914 11104
rect 16945 11101 16957 11104
rect 16991 11101 17003 11135
rect 20548 11132 20576 11163
rect 20714 11160 20720 11212
rect 20772 11160 20778 11212
rect 22094 11160 22100 11212
rect 22152 11160 22158 11212
rect 22370 11160 22376 11212
rect 22428 11160 22434 11212
rect 21174 11132 21180 11144
rect 20548 11104 21180 11132
rect 16945 11095 17003 11101
rect 21174 11092 21180 11104
rect 21232 11092 21238 11144
rect 12989 11067 13047 11073
rect 12989 11033 13001 11067
rect 13035 11064 13047 11067
rect 13722 11064 13728 11076
rect 13035 11036 13728 11064
rect 13035 11033 13047 11036
rect 12989 11027 13047 11033
rect 13722 11024 13728 11036
rect 13780 11024 13786 11076
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 15151 11067 15209 11073
rect 15151 11064 15163 11067
rect 14884 11036 15163 11064
rect 14884 11024 14890 11036
rect 15151 11033 15163 11036
rect 15197 11033 15209 11067
rect 15151 11027 15209 11033
rect 15933 11067 15991 11073
rect 15933 11033 15945 11067
rect 15979 11064 15991 11067
rect 17218 11064 17224 11076
rect 15979 11036 17224 11064
rect 15979 11033 15991 11036
rect 15933 11027 15991 11033
rect 17218 11024 17224 11036
rect 17276 11024 17282 11076
rect 11204 10968 11284 10996
rect 11204 10956 11210 10968
rect 11514 10956 11520 11008
rect 11572 10996 11578 11008
rect 12069 10999 12127 11005
rect 12069 10996 12081 10999
rect 11572 10968 12081 10996
rect 11572 10956 11578 10968
rect 12069 10965 12081 10968
rect 12115 10965 12127 10999
rect 12069 10959 12127 10965
rect 12618 10956 12624 11008
rect 12676 10956 12682 11008
rect 14277 10999 14335 11005
rect 14277 10965 14289 10999
rect 14323 10996 14335 10999
rect 14550 10996 14556 11008
rect 14323 10968 14556 10996
rect 14323 10965 14335 10968
rect 14277 10959 14335 10965
rect 14550 10956 14556 10968
rect 14608 10956 14614 11008
rect 14918 10956 14924 11008
rect 14976 10956 14982 11008
rect 16574 10956 16580 11008
rect 16632 10956 16638 11008
rect 18141 10999 18199 11005
rect 18141 10965 18153 10999
rect 18187 10996 18199 10999
rect 18230 10996 18236 11008
rect 18187 10968 18236 10996
rect 18187 10965 18199 10968
rect 18141 10959 18199 10965
rect 18230 10956 18236 10968
rect 18288 10956 18294 11008
rect 18322 10956 18328 11008
rect 18380 10956 18386 11008
rect 21729 10999 21787 11005
rect 21729 10965 21741 10999
rect 21775 10996 21787 10999
rect 22189 10999 22247 11005
rect 22189 10996 22201 10999
rect 21775 10968 22201 10996
rect 21775 10965 21787 10968
rect 21729 10959 21787 10965
rect 22189 10965 22201 10968
rect 22235 10965 22247 10999
rect 22189 10959 22247 10965
rect 552 10906 23368 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 23368 10906
rect 552 10832 23368 10854
rect 6178 10752 6184 10804
rect 6236 10792 6242 10804
rect 6273 10795 6331 10801
rect 6273 10792 6285 10795
rect 6236 10764 6285 10792
rect 6236 10752 6242 10764
rect 6273 10761 6285 10764
rect 6319 10792 6331 10795
rect 7098 10792 7104 10804
rect 6319 10764 7104 10792
rect 6319 10761 6331 10764
rect 6273 10755 6331 10761
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 9548 10764 9904 10792
rect 9548 10752 9554 10764
rect 4816 10628 5028 10656
rect 3970 10548 3976 10600
rect 4028 10588 4034 10600
rect 4614 10588 4620 10600
rect 4028 10560 4620 10588
rect 4028 10548 4034 10560
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 4816 10597 4844 10628
rect 4801 10591 4859 10597
rect 4801 10557 4813 10591
rect 4847 10557 4859 10591
rect 4801 10551 4859 10557
rect 4246 10480 4252 10532
rect 4304 10520 4310 10532
rect 4816 10520 4844 10551
rect 4890 10548 4896 10600
rect 4948 10548 4954 10600
rect 5000 10588 5028 10628
rect 8294 10616 8300 10668
rect 8352 10656 8358 10668
rect 8481 10659 8539 10665
rect 8481 10656 8493 10659
rect 8352 10628 8493 10656
rect 8352 10616 8358 10628
rect 8481 10625 8493 10628
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 8846 10616 8852 10668
rect 8904 10656 8910 10668
rect 9876 10665 9904 10764
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10502 10792 10508 10804
rect 10008 10764 10508 10792
rect 10008 10752 10014 10764
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 12526 10752 12532 10804
rect 12584 10752 12590 10804
rect 17037 10795 17095 10801
rect 17037 10761 17049 10795
rect 17083 10792 17095 10795
rect 18322 10792 18328 10804
rect 17083 10764 18328 10792
rect 17083 10761 17095 10764
rect 17037 10755 17095 10761
rect 18322 10752 18328 10764
rect 18380 10752 18386 10804
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 21453 10795 21511 10801
rect 21453 10792 21465 10795
rect 20772 10764 21465 10792
rect 20772 10752 20778 10764
rect 21453 10761 21465 10764
rect 21499 10792 21511 10795
rect 22002 10792 22008 10804
rect 21499 10764 22008 10792
rect 21499 10761 21511 10764
rect 21453 10755 21511 10761
rect 22002 10752 22008 10764
rect 22060 10752 22066 10804
rect 22373 10795 22431 10801
rect 22373 10761 22385 10795
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 10410 10684 10416 10736
rect 10468 10684 10474 10736
rect 12391 10727 12449 10733
rect 12391 10724 12403 10727
rect 11808 10696 12403 10724
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 8904 10628 8953 10656
rect 8904 10616 8910 10628
rect 8941 10625 8953 10628
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10656 9919 10659
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 9907 10628 10640 10656
rect 9907 10625 9919 10628
rect 9861 10619 9919 10625
rect 5626 10588 5632 10600
rect 5000 10560 5632 10588
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 6454 10548 6460 10600
rect 6512 10588 6518 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 6512 10560 6561 10588
rect 6512 10548 6518 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8444 10560 8585 10588
rect 8444 10548 8450 10560
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 9766 10588 9772 10600
rect 8573 10551 8631 10557
rect 9324 10560 9772 10588
rect 5166 10529 5172 10532
rect 4304 10492 4844 10520
rect 4304 10480 4310 10492
rect 5160 10483 5172 10529
rect 5166 10480 5172 10483
rect 5224 10480 5230 10532
rect 6362 10480 6368 10532
rect 6420 10480 6426 10532
rect 9324 10529 9352 10560
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10588 10011 10591
rect 10318 10588 10324 10600
rect 9999 10560 10324 10588
rect 9999 10557 10011 10560
rect 9953 10551 10011 10557
rect 10318 10548 10324 10560
rect 10376 10548 10382 10600
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10588 10471 10591
rect 10502 10588 10508 10600
rect 10459 10560 10508 10588
rect 10459 10557 10471 10560
rect 10413 10551 10471 10557
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 10612 10597 10640 10628
rect 11348 10628 11713 10656
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10557 10747 10591
rect 10689 10551 10747 10557
rect 9309 10523 9367 10529
rect 9309 10489 9321 10523
rect 9355 10489 9367 10523
rect 9309 10483 9367 10489
rect 9600 10492 10456 10520
rect 4706 10412 4712 10464
rect 4764 10412 4770 10464
rect 6730 10412 6736 10464
rect 6788 10412 6794 10464
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 9509 10455 9567 10461
rect 9509 10452 9521 10455
rect 9272 10424 9521 10452
rect 9272 10412 9278 10424
rect 9509 10421 9521 10424
rect 9555 10452 9567 10455
rect 9600 10452 9628 10492
rect 9555 10424 9628 10452
rect 9555 10421 9567 10424
rect 9509 10415 9567 10421
rect 9674 10412 9680 10464
rect 9732 10412 9738 10464
rect 10318 10412 10324 10464
rect 10376 10412 10382 10464
rect 10428 10452 10456 10492
rect 10704 10452 10732 10551
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11348 10597 11376 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11333 10591 11391 10597
rect 11333 10588 11345 10591
rect 11112 10560 11345 10588
rect 11112 10548 11118 10560
rect 11333 10557 11345 10560
rect 11379 10557 11391 10591
rect 11333 10551 11391 10557
rect 11514 10548 11520 10600
rect 11572 10548 11578 10600
rect 11808 10597 11836 10696
rect 12391 10693 12403 10696
rect 12437 10724 12449 10727
rect 12618 10724 12624 10736
rect 12437 10696 12624 10724
rect 12437 10693 12449 10696
rect 12391 10687 12449 10693
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 17129 10727 17187 10733
rect 17129 10693 17141 10727
rect 17175 10724 17187 10727
rect 17494 10724 17500 10736
rect 17175 10696 17500 10724
rect 17175 10693 17187 10696
rect 17129 10687 17187 10693
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 14608 10628 15332 10656
rect 14608 10616 14614 10628
rect 11793 10591 11851 10597
rect 11793 10557 11805 10591
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10588 12311 10591
rect 12342 10588 12348 10600
rect 12299 10560 12348 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 12342 10548 12348 10560
rect 12400 10548 12406 10600
rect 12710 10548 12716 10600
rect 12768 10548 12774 10600
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10557 13599 10591
rect 13541 10551 13599 10557
rect 12621 10523 12679 10529
rect 12621 10489 12633 10523
rect 12667 10520 12679 10523
rect 13556 10520 13584 10551
rect 13722 10548 13728 10600
rect 13780 10548 13786 10600
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10588 14703 10591
rect 14826 10588 14832 10600
rect 14691 10560 14832 10588
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 15304 10597 15332 10628
rect 15105 10591 15163 10597
rect 15105 10588 15117 10591
rect 14976 10560 15117 10588
rect 14976 10548 14982 10560
rect 15105 10557 15117 10560
rect 15151 10557 15163 10591
rect 15105 10551 15163 10557
rect 15289 10591 15347 10597
rect 15289 10557 15301 10591
rect 15335 10557 15347 10591
rect 15289 10551 15347 10557
rect 16853 10591 16911 10597
rect 16853 10557 16865 10591
rect 16899 10588 16911 10591
rect 17144 10588 17172 10687
rect 17494 10684 17500 10696
rect 17552 10684 17558 10736
rect 22388 10724 22416 10755
rect 22738 10752 22744 10804
rect 22796 10752 22802 10804
rect 22554 10724 22560 10736
rect 22066 10696 22560 10724
rect 22066 10656 22094 10696
rect 22554 10684 22560 10696
rect 22612 10684 22618 10736
rect 20732 10628 22094 10656
rect 22281 10659 22339 10665
rect 16899 10560 17172 10588
rect 16899 10557 16911 10560
rect 16853 10551 16911 10557
rect 18230 10548 18236 10600
rect 18288 10597 18294 10600
rect 18288 10588 18300 10597
rect 18509 10591 18567 10597
rect 18288 10560 18333 10588
rect 18288 10551 18300 10560
rect 18509 10557 18521 10591
rect 18555 10588 18567 10591
rect 19150 10588 19156 10600
rect 18555 10560 19156 10588
rect 18555 10557 18567 10560
rect 18509 10551 18567 10557
rect 18288 10548 18294 10551
rect 12667 10492 13584 10520
rect 12667 10489 12679 10492
rect 12621 10483 12679 10489
rect 14734 10480 14740 10532
rect 14792 10520 14798 10532
rect 15197 10523 15255 10529
rect 15197 10520 15209 10523
rect 14792 10492 15209 10520
rect 14792 10480 14798 10492
rect 15197 10489 15209 10492
rect 15243 10489 15255 10523
rect 15197 10483 15255 10489
rect 16666 10480 16672 10532
rect 16724 10480 16730 10532
rect 18138 10480 18144 10532
rect 18196 10520 18202 10532
rect 18524 10520 18552 10551
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 18196 10492 18552 10520
rect 20732 10520 20760 10628
rect 22281 10625 22293 10659
rect 22327 10656 22339 10659
rect 22327 10628 22600 10656
rect 22327 10625 22339 10628
rect 22281 10619 22339 10625
rect 20809 10591 20867 10597
rect 20809 10557 20821 10591
rect 20855 10588 20867 10591
rect 21821 10591 21879 10597
rect 20855 10560 21496 10588
rect 20855 10557 20867 10560
rect 20809 10551 20867 10557
rect 20993 10523 21051 10529
rect 20993 10520 21005 10523
rect 20732 10492 21005 10520
rect 18196 10480 18202 10492
rect 20993 10489 21005 10492
rect 21039 10520 21051 10523
rect 21082 10520 21088 10532
rect 21039 10492 21088 10520
rect 21039 10489 21051 10492
rect 20993 10483 21051 10489
rect 21082 10480 21088 10492
rect 21140 10480 21146 10532
rect 21468 10529 21496 10560
rect 21821 10557 21833 10591
rect 21867 10588 21879 10591
rect 21910 10588 21916 10600
rect 21867 10560 21916 10588
rect 21867 10557 21879 10560
rect 21821 10551 21879 10557
rect 21910 10548 21916 10560
rect 21968 10548 21974 10600
rect 22094 10548 22100 10600
rect 22152 10548 22158 10600
rect 22370 10548 22376 10600
rect 22428 10548 22434 10600
rect 22572 10597 22600 10628
rect 22557 10591 22615 10597
rect 22557 10557 22569 10591
rect 22603 10588 22615 10591
rect 22646 10588 22652 10600
rect 22603 10560 22652 10588
rect 22603 10557 22615 10560
rect 22557 10551 22615 10557
rect 22646 10548 22652 10560
rect 22704 10548 22710 10600
rect 21177 10523 21235 10529
rect 21177 10489 21189 10523
rect 21223 10520 21235 10523
rect 21453 10523 21511 10529
rect 21223 10492 21404 10520
rect 21223 10489 21235 10492
rect 21177 10483 21235 10489
rect 10428 10424 10732 10452
rect 11425 10455 11483 10461
rect 11425 10421 11437 10455
rect 11471 10452 11483 10455
rect 11606 10452 11612 10464
rect 11471 10424 11612 10452
rect 11471 10421 11483 10424
rect 11425 10415 11483 10421
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 12158 10412 12164 10464
rect 12216 10412 12222 10464
rect 13722 10412 13728 10464
rect 13780 10412 13786 10464
rect 15013 10455 15071 10461
rect 15013 10421 15025 10455
rect 15059 10452 15071 10455
rect 15102 10452 15108 10464
rect 15059 10424 15108 10452
rect 15059 10421 15071 10424
rect 15013 10415 15071 10421
rect 15102 10412 15108 10424
rect 15160 10412 15166 10464
rect 21266 10412 21272 10464
rect 21324 10412 21330 10464
rect 21376 10452 21404 10492
rect 21453 10489 21465 10523
rect 21499 10489 21511 10523
rect 21453 10483 21511 10489
rect 21913 10455 21971 10461
rect 21913 10452 21925 10455
rect 21376 10424 21925 10452
rect 21913 10421 21925 10424
rect 21959 10452 21971 10455
rect 22462 10452 22468 10464
rect 21959 10424 22468 10452
rect 21959 10421 21971 10424
rect 21913 10415 21971 10421
rect 22462 10412 22468 10424
rect 22520 10412 22526 10464
rect 552 10362 23368 10384
rect 552 10310 4322 10362
rect 4374 10310 4386 10362
rect 4438 10310 4450 10362
rect 4502 10310 4514 10362
rect 4566 10310 4578 10362
rect 4630 10310 23368 10362
rect 552 10288 23368 10310
rect 4341 10251 4399 10257
rect 4341 10217 4353 10251
rect 4387 10248 4399 10251
rect 6362 10248 6368 10260
rect 4387 10220 6368 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 3970 10140 3976 10192
rect 4028 10140 4034 10192
rect 4203 10149 4261 10155
rect 4203 10115 4215 10149
rect 4249 10146 4261 10149
rect 4249 10124 4292 10146
rect 4249 10115 4252 10124
rect 4203 10109 4252 10115
rect 4246 10072 4252 10109
rect 4304 10072 4310 10124
rect 4448 10121 4476 10220
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 9861 10251 9919 10257
rect 9861 10217 9873 10251
rect 9907 10248 9919 10251
rect 9907 10220 12204 10248
rect 9907 10217 9919 10220
rect 9861 10211 9919 10217
rect 4798 10140 4804 10192
rect 4856 10140 4862 10192
rect 5074 10140 5080 10192
rect 5132 10140 5138 10192
rect 5353 10183 5411 10189
rect 5353 10149 5365 10183
rect 5399 10180 5411 10183
rect 5399 10152 5948 10180
rect 5399 10149 5411 10152
rect 5353 10143 5411 10149
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10081 4491 10115
rect 5258 10112 5264 10124
rect 4433 10075 4491 10081
rect 4724 10084 5264 10112
rect 4724 10044 4752 10084
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5368 10084 5457 10112
rect 5368 10056 5396 10084
rect 5445 10081 5457 10084
rect 5491 10112 5503 10115
rect 5626 10112 5632 10124
rect 5491 10084 5632 10112
rect 5491 10081 5503 10084
rect 5445 10075 5503 10081
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 4172 10016 4752 10044
rect 4172 9917 4200 10016
rect 5350 10004 5356 10056
rect 5408 10004 5414 10056
rect 5810 10004 5816 10056
rect 5868 10004 5874 10056
rect 5828 9976 5856 10004
rect 4816 9948 5856 9976
rect 4816 9917 4844 9948
rect 4157 9911 4215 9917
rect 4157 9877 4169 9911
rect 4203 9877 4215 9911
rect 4157 9871 4215 9877
rect 4801 9911 4859 9917
rect 4801 9877 4813 9911
rect 4847 9877 4859 9911
rect 4801 9871 4859 9877
rect 4982 9868 4988 9920
rect 5040 9868 5046 9920
rect 5626 9868 5632 9920
rect 5684 9868 5690 9920
rect 5813 9911 5871 9917
rect 5813 9877 5825 9911
rect 5859 9908 5871 9911
rect 5920 9908 5948 10152
rect 9306 10140 9312 10192
rect 9364 10180 9370 10192
rect 12176 10189 12204 10220
rect 16390 10208 16396 10260
rect 16448 10208 16454 10260
rect 16853 10251 16911 10257
rect 16853 10217 16865 10251
rect 16899 10248 16911 10251
rect 17034 10248 17040 10260
rect 16899 10220 17040 10248
rect 16899 10217 16911 10220
rect 16853 10211 16911 10217
rect 9401 10183 9459 10189
rect 9401 10180 9413 10183
rect 9364 10152 9413 10180
rect 9364 10140 9370 10152
rect 9401 10149 9413 10152
rect 9447 10149 9459 10183
rect 9401 10143 9459 10149
rect 12161 10183 12219 10189
rect 12161 10149 12173 10183
rect 12207 10149 12219 10183
rect 12161 10143 12219 10149
rect 6914 10072 6920 10124
rect 6972 10121 6978 10124
rect 6972 10075 6984 10121
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10112 7251 10115
rect 8662 10112 8668 10124
rect 7239 10084 8668 10112
rect 7239 10081 7251 10084
rect 7193 10075 7251 10081
rect 6972 10072 6978 10075
rect 8662 10072 8668 10084
rect 8720 10072 8726 10124
rect 8754 10072 8760 10124
rect 8812 10072 8818 10124
rect 9674 10072 9680 10124
rect 9732 10072 9738 10124
rect 11698 10072 11704 10124
rect 11756 10072 11762 10124
rect 12434 10072 12440 10124
rect 12492 10072 12498 10124
rect 13814 10072 13820 10124
rect 13872 10072 13878 10124
rect 14550 10072 14556 10124
rect 14608 10072 14614 10124
rect 15197 10115 15255 10121
rect 15197 10081 15209 10115
rect 15243 10112 15255 10115
rect 15378 10112 15384 10124
rect 15243 10084 15384 10112
rect 15243 10081 15255 10084
rect 15197 10075 15255 10081
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 16298 10072 16304 10124
rect 16356 10072 16362 10124
rect 16577 10115 16635 10121
rect 16577 10081 16589 10115
rect 16623 10112 16635 10115
rect 16868 10112 16896 10211
rect 17034 10208 17040 10220
rect 17092 10248 17098 10260
rect 17770 10248 17776 10260
rect 17092 10220 17776 10248
rect 17092 10208 17098 10220
rect 17770 10208 17776 10220
rect 17828 10208 17834 10260
rect 21269 10251 21327 10257
rect 21269 10217 21281 10251
rect 21315 10248 21327 10251
rect 21450 10248 21456 10260
rect 21315 10220 21456 10248
rect 21315 10217 21327 10220
rect 21269 10211 21327 10217
rect 21450 10208 21456 10220
rect 21508 10208 21514 10260
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 22097 10251 22155 10257
rect 22097 10248 22109 10251
rect 22060 10220 22109 10248
rect 22060 10208 22066 10220
rect 22097 10217 22109 10220
rect 22143 10217 22155 10251
rect 22097 10211 22155 10217
rect 22186 10208 22192 10260
rect 22244 10248 22250 10260
rect 22244 10220 22600 10248
rect 22244 10208 22250 10220
rect 21082 10140 21088 10192
rect 21140 10140 21146 10192
rect 22572 10189 22600 10220
rect 22557 10183 22615 10189
rect 22557 10149 22569 10183
rect 22603 10149 22615 10183
rect 22557 10143 22615 10149
rect 16623 10084 16896 10112
rect 16623 10081 16635 10084
rect 16577 10075 16635 10081
rect 17494 10072 17500 10124
rect 17552 10112 17558 10124
rect 17966 10115 18024 10121
rect 17966 10112 17978 10115
rect 17552 10084 17978 10112
rect 17552 10072 17558 10084
rect 17966 10081 17978 10084
rect 18012 10081 18024 10115
rect 17966 10075 18024 10081
rect 18138 10072 18144 10124
rect 18196 10112 18202 10124
rect 18233 10115 18291 10121
rect 18233 10112 18245 10115
rect 18196 10084 18245 10112
rect 18196 10072 18202 10084
rect 18233 10081 18245 10084
rect 18279 10081 18291 10115
rect 18233 10075 18291 10081
rect 19705 10115 19763 10121
rect 19705 10081 19717 10115
rect 19751 10112 19763 10115
rect 20254 10112 20260 10124
rect 19751 10084 20260 10112
rect 19751 10081 19763 10084
rect 19705 10075 19763 10081
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 20717 10115 20775 10121
rect 20717 10112 20729 10115
rect 20456 10084 20729 10112
rect 8846 10004 8852 10056
rect 8904 10004 8910 10056
rect 9493 10047 9551 10053
rect 9493 10044 9505 10047
rect 9140 10016 9505 10044
rect 9140 9985 9168 10016
rect 9493 10013 9505 10016
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 11606 10004 11612 10056
rect 11664 10004 11670 10056
rect 12250 10004 12256 10056
rect 12308 10004 12314 10056
rect 13722 10004 13728 10056
rect 13780 10004 13786 10056
rect 14645 10047 14703 10053
rect 14645 10013 14657 10047
rect 14691 10044 14703 10047
rect 14734 10044 14740 10056
rect 14691 10016 14740 10044
rect 14691 10013 14703 10016
rect 14645 10007 14703 10013
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 15102 10004 15108 10056
rect 15160 10004 15166 10056
rect 19886 10004 19892 10056
rect 19944 10044 19950 10056
rect 20456 10044 20484 10084
rect 20717 10081 20729 10084
rect 20763 10081 20775 10115
rect 20717 10075 20775 10081
rect 20806 10072 20812 10124
rect 20864 10072 20870 10124
rect 20898 10072 20904 10124
rect 20956 10072 20962 10124
rect 21637 10115 21695 10121
rect 21637 10081 21649 10115
rect 21683 10112 21695 10115
rect 21683 10084 22416 10112
rect 21683 10081 21695 10084
rect 21637 10075 21695 10081
rect 19944 10016 20484 10044
rect 20533 10047 20591 10053
rect 19944 10004 19950 10016
rect 20533 10013 20545 10047
rect 20579 10044 20591 10047
rect 21453 10047 21511 10053
rect 21453 10044 21465 10047
rect 20579 10016 21465 10044
rect 20579 10013 20591 10016
rect 20533 10007 20591 10013
rect 21453 10013 21465 10016
rect 21499 10013 21511 10047
rect 21453 10007 21511 10013
rect 21542 10004 21548 10056
rect 21600 10004 21606 10056
rect 21729 10047 21787 10053
rect 21729 10013 21741 10047
rect 21775 10044 21787 10047
rect 22388 10044 22416 10084
rect 22462 10072 22468 10124
rect 22520 10072 22526 10124
rect 22646 10072 22652 10124
rect 22704 10112 22710 10124
rect 22741 10115 22799 10121
rect 22741 10112 22753 10115
rect 22704 10084 22753 10112
rect 22704 10072 22710 10084
rect 22741 10081 22753 10084
rect 22787 10081 22799 10115
rect 22741 10075 22799 10081
rect 22664 10044 22692 10072
rect 21775 10016 22094 10044
rect 22388 10016 22692 10044
rect 21775 10013 21787 10016
rect 21729 10007 21787 10013
rect 9125 9979 9183 9985
rect 9125 9945 9137 9979
rect 9171 9945 9183 9979
rect 9125 9939 9183 9945
rect 14185 9979 14243 9985
rect 14185 9945 14197 9979
rect 14231 9976 14243 9979
rect 15194 9976 15200 9988
rect 14231 9948 15200 9976
rect 14231 9945 14243 9948
rect 14185 9939 14243 9945
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 22066 9976 22094 10016
rect 22830 9976 22836 9988
rect 22066 9948 22836 9976
rect 22830 9936 22836 9948
rect 22888 9936 22894 9988
rect 6454 9908 6460 9920
rect 5859 9880 6460 9908
rect 5859 9877 5871 9880
rect 5813 9871 5871 9877
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 9677 9911 9735 9917
rect 9677 9877 9689 9911
rect 9723 9908 9735 9911
rect 10410 9908 10416 9920
rect 9723 9880 10416 9908
rect 9723 9877 9735 9880
rect 9677 9871 9735 9877
rect 10410 9868 10416 9880
rect 10468 9868 10474 9920
rect 11977 9911 12035 9917
rect 11977 9877 11989 9911
rect 12023 9908 12035 9911
rect 12161 9911 12219 9917
rect 12161 9908 12173 9911
rect 12023 9880 12173 9908
rect 12023 9877 12035 9880
rect 11977 9871 12035 9877
rect 12161 9877 12173 9880
rect 12207 9877 12219 9911
rect 12161 9871 12219 9877
rect 12621 9911 12679 9917
rect 12621 9877 12633 9911
rect 12667 9908 12679 9911
rect 14734 9908 14740 9920
rect 12667 9880 14740 9908
rect 12667 9877 12679 9880
rect 12621 9871 12679 9877
rect 14734 9868 14740 9880
rect 14792 9868 14798 9920
rect 14826 9868 14832 9920
rect 14884 9868 14890 9920
rect 15286 9868 15292 9920
rect 15344 9908 15350 9920
rect 15473 9911 15531 9917
rect 15473 9908 15485 9911
rect 15344 9880 15485 9908
rect 15344 9868 15350 9880
rect 15473 9877 15485 9880
rect 15519 9877 15531 9911
rect 15473 9871 15531 9877
rect 16758 9868 16764 9920
rect 16816 9868 16822 9920
rect 19521 9911 19579 9917
rect 19521 9877 19533 9911
rect 19567 9908 19579 9911
rect 19610 9908 19616 9920
rect 19567 9880 19616 9908
rect 19567 9877 19579 9880
rect 19521 9871 19579 9877
rect 19610 9868 19616 9880
rect 19668 9868 19674 9920
rect 21818 9868 21824 9920
rect 21876 9908 21882 9920
rect 21913 9911 21971 9917
rect 21913 9908 21925 9911
rect 21876 9880 21925 9908
rect 21876 9868 21882 9880
rect 21913 9877 21925 9880
rect 21959 9877 21971 9911
rect 21913 9871 21971 9877
rect 22097 9911 22155 9917
rect 22097 9877 22109 9911
rect 22143 9908 22155 9911
rect 22925 9911 22983 9917
rect 22925 9908 22937 9911
rect 22143 9880 22937 9908
rect 22143 9877 22155 9880
rect 22097 9871 22155 9877
rect 22925 9877 22937 9880
rect 22971 9877 22983 9911
rect 22925 9871 22983 9877
rect 552 9818 23368 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 23368 9818
rect 552 9744 23368 9766
rect 4617 9707 4675 9713
rect 4617 9673 4629 9707
rect 4663 9704 4675 9707
rect 4706 9704 4712 9716
rect 4663 9676 4712 9704
rect 4663 9673 4675 9676
rect 4617 9667 4675 9673
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 4801 9707 4859 9713
rect 4801 9673 4813 9707
rect 4847 9704 4859 9707
rect 5166 9704 5172 9716
rect 4847 9676 5172 9704
rect 4847 9673 4859 9676
rect 4801 9667 4859 9673
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 5994 9704 6000 9716
rect 5316 9676 6000 9704
rect 5316 9664 5322 9676
rect 5994 9664 6000 9676
rect 6052 9704 6058 9716
rect 6052 9676 6316 9704
rect 6052 9664 6058 9676
rect 6288 9645 6316 9676
rect 6730 9664 6736 9716
rect 6788 9664 6794 9716
rect 6914 9664 6920 9716
rect 6972 9664 6978 9716
rect 8757 9707 8815 9713
rect 8757 9673 8769 9707
rect 8803 9704 8815 9707
rect 9950 9704 9956 9716
rect 8803 9676 9956 9704
rect 8803 9673 8815 9676
rect 8757 9667 8815 9673
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 11333 9707 11391 9713
rect 11333 9673 11345 9707
rect 11379 9704 11391 9707
rect 12250 9704 12256 9716
rect 11379 9676 12256 9704
rect 11379 9673 11391 9676
rect 11333 9667 11391 9673
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 14369 9707 14427 9713
rect 14369 9673 14381 9707
rect 14415 9704 14427 9707
rect 14642 9704 14648 9716
rect 14415 9676 14648 9704
rect 14415 9673 14427 9676
rect 14369 9667 14427 9673
rect 14642 9664 14648 9676
rect 14700 9664 14706 9716
rect 14826 9664 14832 9716
rect 14884 9704 14890 9716
rect 15013 9707 15071 9713
rect 15013 9704 15025 9707
rect 14884 9676 15025 9704
rect 14884 9664 14890 9676
rect 15013 9673 15025 9676
rect 15059 9673 15071 9707
rect 15013 9667 15071 9673
rect 16758 9664 16764 9716
rect 16816 9704 16822 9716
rect 17313 9707 17371 9713
rect 17313 9704 17325 9707
rect 16816 9676 17325 9704
rect 16816 9664 16822 9676
rect 17313 9673 17325 9676
rect 17359 9673 17371 9707
rect 17589 9707 17647 9713
rect 17589 9704 17601 9707
rect 17313 9667 17371 9673
rect 17420 9676 17601 9704
rect 6273 9639 6331 9645
rect 6273 9605 6285 9639
rect 6319 9605 6331 9639
rect 6273 9599 6331 9605
rect 12434 9596 12440 9648
rect 12492 9596 12498 9648
rect 14458 9596 14464 9648
rect 14516 9636 14522 9648
rect 14553 9639 14611 9645
rect 14553 9636 14565 9639
rect 14516 9608 14565 9636
rect 14516 9596 14522 9608
rect 14553 9605 14565 9608
rect 14599 9605 14611 9639
rect 14553 9599 14611 9605
rect 15473 9639 15531 9645
rect 15473 9605 15485 9639
rect 15519 9636 15531 9639
rect 16574 9636 16580 9648
rect 15519 9608 16580 9636
rect 15519 9605 15531 9608
rect 15473 9599 15531 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 16945 9639 17003 9645
rect 16945 9636 16957 9639
rect 16724 9608 16957 9636
rect 16724 9596 16730 9608
rect 16945 9605 16957 9608
rect 16991 9636 17003 9639
rect 17420 9636 17448 9676
rect 17589 9673 17601 9676
rect 17635 9673 17647 9707
rect 17589 9667 17647 9673
rect 17770 9664 17776 9716
rect 17828 9664 17834 9716
rect 18230 9664 18236 9716
rect 18288 9704 18294 9716
rect 18414 9704 18420 9716
rect 18288 9676 18420 9704
rect 18288 9664 18294 9676
rect 18414 9664 18420 9676
rect 18472 9704 18478 9716
rect 19242 9704 19248 9716
rect 18472 9676 19248 9704
rect 18472 9664 18478 9676
rect 19242 9664 19248 9676
rect 19300 9664 19306 9716
rect 19812 9676 20760 9704
rect 16991 9608 17448 9636
rect 16991 9605 17003 9608
rect 16945 9599 17003 9605
rect 17494 9596 17500 9648
rect 17552 9596 17558 9648
rect 4890 9528 4896 9580
rect 4948 9528 4954 9580
rect 10318 9528 10324 9580
rect 10376 9568 10382 9580
rect 10873 9571 10931 9577
rect 10873 9568 10885 9571
rect 10376 9540 10885 9568
rect 10376 9528 10382 9540
rect 10873 9537 10885 9540
rect 10919 9537 10931 9571
rect 10873 9531 10931 9537
rect 12158 9528 12164 9580
rect 12216 9528 12222 9580
rect 15194 9528 15200 9580
rect 15252 9528 15258 9580
rect 16390 9528 16396 9580
rect 16448 9568 16454 9580
rect 16448 9540 16896 9568
rect 16448 9528 16454 9540
rect 4982 9460 4988 9512
rect 5040 9500 5046 9512
rect 5149 9503 5207 9509
rect 5149 9500 5161 9503
rect 5040 9472 5161 9500
rect 5040 9460 5046 9472
rect 5149 9469 5161 9472
rect 5195 9469 5207 9503
rect 5149 9463 5207 9469
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 5684 9472 6377 9500
rect 5684 9460 5690 9472
rect 6365 9469 6377 9472
rect 6411 9500 6423 9503
rect 7650 9500 7656 9512
rect 6411 9472 7656 9500
rect 6411 9469 6423 9472
rect 6365 9463 6423 9469
rect 7650 9460 7656 9472
rect 7708 9500 7714 9512
rect 7929 9503 7987 9509
rect 7929 9500 7941 9503
rect 7708 9472 7941 9500
rect 7708 9460 7714 9472
rect 7929 9469 7941 9472
rect 7975 9469 7987 9503
rect 7929 9463 7987 9469
rect 8386 9460 8392 9512
rect 8444 9500 8450 9512
rect 9033 9503 9091 9509
rect 9033 9500 9045 9503
rect 8444 9472 9045 9500
rect 8444 9460 8450 9472
rect 9033 9469 9045 9472
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9766 9500 9772 9512
rect 9263 9472 9772 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10888 9472 10977 9500
rect 10888 9444 10916 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 12066 9460 12072 9512
rect 12124 9460 12130 9512
rect 14734 9460 14740 9512
rect 14792 9500 14798 9512
rect 15013 9503 15071 9509
rect 15013 9500 15025 9503
rect 14792 9472 15025 9500
rect 14792 9460 14798 9472
rect 15013 9469 15025 9472
rect 15059 9469 15071 9503
rect 15013 9463 15071 9469
rect 15286 9460 15292 9512
rect 15344 9460 15350 9512
rect 15470 9460 15476 9512
rect 15528 9500 15534 9512
rect 16298 9500 16304 9512
rect 15528 9472 16304 9500
rect 15528 9460 15534 9472
rect 16298 9460 16304 9472
rect 16356 9500 16362 9512
rect 16482 9500 16488 9512
rect 16356 9472 16488 9500
rect 16356 9460 16362 9472
rect 16482 9460 16488 9472
rect 16540 9500 16546 9512
rect 16868 9509 16896 9540
rect 17034 9528 17040 9580
rect 17092 9568 17098 9580
rect 19812 9568 19840 9676
rect 20732 9636 20760 9676
rect 20806 9664 20812 9716
rect 20864 9704 20870 9716
rect 21177 9707 21235 9713
rect 21177 9704 21189 9707
rect 20864 9676 21189 9704
rect 20864 9664 20870 9676
rect 21177 9673 21189 9676
rect 21223 9673 21235 9707
rect 21177 9667 21235 9673
rect 20990 9636 20996 9648
rect 20732 9608 20996 9636
rect 20990 9596 20996 9608
rect 21048 9596 21054 9648
rect 17092 9540 19840 9568
rect 17092 9528 17098 9540
rect 16669 9503 16727 9509
rect 16669 9500 16681 9503
rect 16540 9472 16681 9500
rect 16540 9460 16546 9472
rect 16669 9469 16681 9472
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 16853 9503 16911 9509
rect 16853 9469 16865 9503
rect 16899 9500 16911 9503
rect 18785 9503 18843 9509
rect 16899 9472 18000 9500
rect 16899 9469 16911 9472
rect 16853 9463 16911 9469
rect 4433 9435 4491 9441
rect 4433 9401 4445 9435
rect 4479 9401 4491 9435
rect 4433 9395 4491 9401
rect 4649 9435 4707 9441
rect 4649 9401 4661 9435
rect 4695 9432 4707 9435
rect 5258 9432 5264 9444
rect 4695 9404 5264 9432
rect 4695 9401 4707 9404
rect 4649 9395 4707 9401
rect 4448 9364 4476 9395
rect 5258 9392 5264 9404
rect 5316 9392 5322 9444
rect 6733 9435 6791 9441
rect 6733 9401 6745 9435
rect 6779 9432 6791 9435
rect 6914 9432 6920 9444
rect 6779 9404 6920 9432
rect 6779 9401 6791 9404
rect 6733 9395 6791 9401
rect 6914 9392 6920 9404
rect 6972 9432 6978 9444
rect 7745 9435 7803 9441
rect 6972 9404 7696 9432
rect 6972 9392 6978 9404
rect 4798 9364 4804 9376
rect 4448 9336 4804 9364
rect 4798 9324 4804 9336
rect 4856 9364 4862 9376
rect 5166 9364 5172 9376
rect 4856 9336 5172 9364
rect 4856 9324 4862 9336
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 7558 9324 7564 9376
rect 7616 9324 7622 9376
rect 7668 9364 7696 9404
rect 7745 9401 7757 9435
rect 7791 9432 7803 9435
rect 8570 9432 8576 9444
rect 7791 9404 8576 9432
rect 7791 9401 7803 9404
rect 7745 9395 7803 9401
rect 8570 9392 8576 9404
rect 8628 9392 8634 9444
rect 10870 9392 10876 9444
rect 10928 9392 10934 9444
rect 13814 9392 13820 9444
rect 13872 9432 13878 9444
rect 14185 9435 14243 9441
rect 14185 9432 14197 9435
rect 13872 9404 14197 9432
rect 13872 9392 13878 9404
rect 14185 9401 14197 9404
rect 14231 9401 14243 9435
rect 14185 9395 14243 9401
rect 14274 9392 14280 9444
rect 14332 9432 14338 9444
rect 14401 9435 14459 9441
rect 14401 9432 14413 9435
rect 14332 9404 14413 9432
rect 14332 9392 14338 9404
rect 14401 9401 14413 9404
rect 14447 9432 14459 9435
rect 14918 9432 14924 9444
rect 14447 9404 14924 9432
rect 14447 9401 14459 9404
rect 14401 9395 14459 9401
rect 14918 9392 14924 9404
rect 14976 9392 14982 9444
rect 16684 9432 16712 9463
rect 17757 9435 17815 9441
rect 17757 9432 17769 9435
rect 16684 9404 17769 9432
rect 17757 9401 17769 9404
rect 17803 9432 17815 9435
rect 17862 9432 17868 9444
rect 17803 9404 17868 9432
rect 17803 9401 17815 9404
rect 17757 9395 17815 9401
rect 17862 9392 17868 9404
rect 17920 9392 17926 9444
rect 17972 9441 18000 9472
rect 18785 9469 18797 9503
rect 18831 9469 18843 9503
rect 18785 9463 18843 9469
rect 18969 9503 19027 9509
rect 18969 9469 18981 9503
rect 19015 9500 19027 9503
rect 19610 9500 19616 9512
rect 19015 9472 19616 9500
rect 19015 9469 19027 9472
rect 18969 9463 19027 9469
rect 17957 9435 18015 9441
rect 17957 9401 17969 9435
rect 18003 9401 18015 9435
rect 18800 9432 18828 9463
rect 19610 9460 19616 9472
rect 19668 9460 19674 9512
rect 19797 9503 19855 9509
rect 19797 9469 19809 9503
rect 19843 9500 19855 9503
rect 19884 9500 20024 9502
rect 21174 9500 21180 9512
rect 19843 9474 21180 9500
rect 19843 9472 19912 9474
rect 19996 9472 21180 9474
rect 19843 9469 19855 9472
rect 19797 9463 19855 9469
rect 21174 9460 21180 9472
rect 21232 9500 21238 9512
rect 21818 9509 21824 9512
rect 21545 9503 21603 9509
rect 21545 9500 21557 9503
rect 21232 9472 21557 9500
rect 21232 9460 21238 9472
rect 21545 9469 21557 9472
rect 21591 9469 21603 9503
rect 21812 9500 21824 9509
rect 21779 9472 21824 9500
rect 21545 9463 21603 9469
rect 21812 9463 21824 9472
rect 21818 9460 21824 9463
rect 21876 9460 21882 9512
rect 20064 9435 20122 9441
rect 18800 9404 19840 9432
rect 17957 9395 18015 9401
rect 19812 9376 19840 9404
rect 20064 9401 20076 9435
rect 20110 9432 20122 9435
rect 20162 9432 20168 9444
rect 20110 9404 20168 9432
rect 20110 9401 20122 9404
rect 20064 9395 20122 9401
rect 20162 9392 20168 9404
rect 20220 9392 20226 9444
rect 8202 9364 8208 9376
rect 7668 9336 8208 9364
rect 8202 9324 8208 9336
rect 8260 9364 8266 9376
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 8260 9336 8769 9364
rect 8260 9324 8266 9336
rect 8757 9333 8769 9336
rect 8803 9333 8815 9367
rect 8757 9327 8815 9333
rect 8938 9324 8944 9376
rect 8996 9324 9002 9376
rect 9401 9367 9459 9373
rect 9401 9333 9413 9367
rect 9447 9364 9459 9367
rect 9490 9364 9496 9376
rect 9447 9336 9496 9364
rect 9447 9333 9459 9336
rect 9401 9327 9459 9333
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 12986 9324 12992 9376
rect 13044 9364 13050 9376
rect 16758 9364 16764 9376
rect 13044 9336 16764 9364
rect 13044 9324 13050 9336
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 16850 9324 16856 9376
rect 16908 9324 16914 9376
rect 17310 9324 17316 9376
rect 17368 9324 17374 9376
rect 18782 9324 18788 9376
rect 18840 9324 18846 9376
rect 19061 9367 19119 9373
rect 19061 9333 19073 9367
rect 19107 9364 19119 9367
rect 19150 9364 19156 9376
rect 19107 9336 19156 9364
rect 19107 9333 19119 9336
rect 19061 9327 19119 9333
rect 19150 9324 19156 9336
rect 19208 9324 19214 9376
rect 19245 9367 19303 9373
rect 19245 9333 19257 9367
rect 19291 9364 19303 9367
rect 19702 9364 19708 9376
rect 19291 9336 19708 9364
rect 19291 9333 19303 9336
rect 19245 9327 19303 9333
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 19794 9324 19800 9376
rect 19852 9324 19858 9376
rect 19978 9324 19984 9376
rect 20036 9364 20042 9376
rect 20530 9364 20536 9376
rect 20036 9336 20536 9364
rect 20036 9324 20042 9336
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 22646 9324 22652 9376
rect 22704 9364 22710 9376
rect 22925 9367 22983 9373
rect 22925 9364 22937 9367
rect 22704 9336 22937 9364
rect 22704 9324 22710 9336
rect 22925 9333 22937 9336
rect 22971 9333 22983 9367
rect 22925 9327 22983 9333
rect 552 9274 23368 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 23368 9274
rect 552 9200 23368 9222
rect 5258 9120 5264 9172
rect 5316 9120 5322 9172
rect 7127 9163 7185 9169
rect 7127 9129 7139 9163
rect 7173 9160 7185 9163
rect 7558 9160 7564 9172
rect 7173 9132 7564 9160
rect 7173 9129 7185 9132
rect 7127 9123 7185 9129
rect 7558 9120 7564 9132
rect 7616 9120 7622 9172
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9766 9160 9772 9172
rect 9171 9132 9772 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 9950 9120 9956 9172
rect 10008 9120 10014 9172
rect 10778 9160 10784 9172
rect 10152 9132 10784 9160
rect 5074 9052 5080 9104
rect 5132 9092 5138 9104
rect 5445 9095 5503 9101
rect 5445 9092 5457 9095
rect 5132 9064 5457 9092
rect 5132 9052 5138 9064
rect 5445 9061 5457 9064
rect 5491 9061 5503 9095
rect 6914 9092 6920 9104
rect 5445 9055 5503 9061
rect 5736 9064 6920 9092
rect 5350 8984 5356 9036
rect 5408 9024 5414 9036
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 5408 8996 5641 9024
rect 5408 8984 5414 8996
rect 5629 8993 5641 8996
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 5736 8956 5764 9064
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 7742 9052 7748 9104
rect 7800 9052 7806 9104
rect 7834 9052 7840 9104
rect 7892 9092 7898 9104
rect 8754 9092 8760 9104
rect 7892 9064 8760 9092
rect 7892 9052 7898 9064
rect 8754 9052 8760 9064
rect 8812 9092 8818 9104
rect 9033 9095 9091 9101
rect 9033 9092 9045 9095
rect 8812 9064 9045 9092
rect 8812 9052 8818 9064
rect 9033 9061 9045 9064
rect 9079 9092 9091 9095
rect 9079 9064 9812 9092
rect 9079 9061 9091 9064
rect 9033 9055 9091 9061
rect 7633 9027 7691 9033
rect 7633 9024 7645 9027
rect 5316 8928 5764 8956
rect 7300 8996 7645 9024
rect 5316 8916 5322 8928
rect 7300 8897 7328 8996
rect 7633 8993 7645 8996
rect 7679 8993 7691 9027
rect 7760 9024 7788 9052
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 7760 8996 9229 9024
rect 7633 8987 7691 8993
rect 9217 8993 9229 8996
rect 9263 9024 9275 9027
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 9263 8996 9505 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 9582 8984 9588 9036
rect 9640 8984 9646 9036
rect 9784 9033 9812 9064
rect 10152 9033 10180 9132
rect 10778 9120 10784 9132
rect 10836 9160 10842 9172
rect 11133 9163 11191 9169
rect 11133 9160 11145 9163
rect 10836 9132 11145 9160
rect 10836 9120 10842 9132
rect 11133 9129 11145 9132
rect 11179 9160 11191 9163
rect 11793 9163 11851 9169
rect 11793 9160 11805 9163
rect 11179 9132 11805 9160
rect 11179 9129 11191 9132
rect 11133 9123 11191 9129
rect 11793 9129 11805 9132
rect 11839 9129 11851 9163
rect 11793 9123 11851 9129
rect 12066 9120 12072 9172
rect 12124 9120 12130 9172
rect 18443 9163 18501 9169
rect 13280 9132 18368 9160
rect 10597 9095 10655 9101
rect 10597 9061 10609 9095
rect 10643 9092 10655 9095
rect 11333 9095 11391 9101
rect 10643 9064 10916 9092
rect 10643 9061 10655 9064
rect 10597 9055 10655 9061
rect 9769 9027 9827 9033
rect 9769 8993 9781 9027
rect 9815 8993 9827 9027
rect 9769 8987 9827 8993
rect 10137 9027 10195 9033
rect 10137 8993 10149 9027
rect 10183 8993 10195 9027
rect 10137 8987 10195 8993
rect 10321 9027 10379 9033
rect 10321 8993 10333 9027
rect 10367 9024 10379 9027
rect 10612 9024 10640 9055
rect 10888 9036 10916 9064
rect 11333 9061 11345 9095
rect 11379 9092 11391 9095
rect 11701 9095 11759 9101
rect 11379 9064 11413 9092
rect 11379 9061 11391 9064
rect 11333 9055 11391 9061
rect 11701 9061 11713 9095
rect 11747 9092 11759 9095
rect 12084 9092 12112 9120
rect 11747 9064 12296 9092
rect 11747 9061 11759 9064
rect 11701 9055 11759 9061
rect 10367 8996 10640 9024
rect 10367 8993 10379 8996
rect 10321 8987 10379 8993
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 10152 8956 10180 8987
rect 10778 8984 10784 9036
rect 10836 8984 10842 9036
rect 10870 8984 10876 9036
rect 10928 9024 10934 9036
rect 11348 9024 11376 9055
rect 11425 9027 11483 9033
rect 11425 9024 11437 9027
rect 10928 8996 11437 9024
rect 10928 8984 10934 8996
rect 11425 8993 11437 8996
rect 11471 8993 11483 9027
rect 11425 8987 11483 8993
rect 11606 8984 11612 9036
rect 11664 8984 11670 9036
rect 12268 9033 12296 9064
rect 13078 9052 13084 9104
rect 13136 9052 13142 9104
rect 13280 9101 13308 9132
rect 13265 9095 13323 9101
rect 13265 9061 13277 9095
rect 13311 9061 13323 9095
rect 14093 9095 14151 9101
rect 13265 9055 13323 9061
rect 13556 9064 13860 9092
rect 12069 9027 12127 9033
rect 12069 8993 12081 9027
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 12253 9027 12311 9033
rect 12253 8993 12265 9027
rect 12299 9024 12311 9027
rect 12802 9024 12808 9036
rect 12299 8996 12808 9024
rect 12299 8993 12311 8996
rect 12253 8987 12311 8993
rect 12084 8956 12112 8987
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 9447 8928 10180 8956
rect 10980 8928 12112 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 7285 8891 7343 8897
rect 7285 8857 7297 8891
rect 7331 8857 7343 8891
rect 7285 8851 7343 8857
rect 7098 8780 7104 8832
rect 7156 8780 7162 8832
rect 7392 8820 7420 8919
rect 8570 8848 8576 8900
rect 8628 8888 8634 8900
rect 8757 8891 8815 8897
rect 8757 8888 8769 8891
rect 8628 8860 8769 8888
rect 8628 8848 8634 8860
rect 8757 8857 8769 8860
rect 8803 8888 8815 8891
rect 8849 8891 8907 8897
rect 8849 8888 8861 8891
rect 8803 8860 8861 8888
rect 8803 8857 8815 8860
rect 8757 8851 8815 8857
rect 8849 8857 8861 8860
rect 8895 8888 8907 8891
rect 9582 8888 9588 8900
rect 8895 8860 9588 8888
rect 8895 8857 8907 8860
rect 8849 8851 8907 8857
rect 9582 8848 9588 8860
rect 9640 8848 9646 8900
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 10980 8897 11008 8928
rect 10965 8891 11023 8897
rect 10965 8888 10977 8891
rect 10744 8860 10977 8888
rect 10744 8848 10750 8860
rect 10965 8857 10977 8860
rect 11011 8857 11023 8891
rect 11606 8888 11612 8900
rect 10965 8851 11023 8857
rect 11164 8860 11612 8888
rect 8662 8820 8668 8832
rect 7392 8792 8668 8820
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 10226 8780 10232 8832
rect 10284 8780 10290 8832
rect 10413 8823 10471 8829
rect 10413 8789 10425 8823
rect 10459 8820 10471 8823
rect 10594 8820 10600 8832
rect 10459 8792 10600 8820
rect 10459 8789 10471 8792
rect 10413 8783 10471 8789
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 11164 8829 11192 8860
rect 11606 8848 11612 8860
rect 11664 8848 11670 8900
rect 13556 8888 13584 9064
rect 13633 9027 13691 9033
rect 13633 8993 13645 9027
rect 13679 9024 13691 9027
rect 13722 9024 13728 9036
rect 13679 8996 13728 9024
rect 13679 8993 13691 8996
rect 13633 8987 13691 8993
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 13832 9033 13860 9064
rect 14093 9061 14105 9095
rect 14139 9092 14151 9095
rect 15197 9095 15255 9101
rect 15197 9092 15209 9095
rect 14139 9064 14412 9092
rect 14139 9061 14151 9064
rect 14093 9055 14151 9061
rect 13817 9027 13875 9033
rect 13817 8993 13829 9027
rect 13863 9024 13875 9027
rect 14274 9024 14280 9036
rect 13863 8996 14280 9024
rect 13863 8993 13875 8996
rect 13817 8987 13875 8993
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 11992 8860 13584 8888
rect 13740 8888 13768 8984
rect 14384 8956 14412 9064
rect 14476 9064 15209 9092
rect 14476 9036 14504 9064
rect 15197 9061 15209 9064
rect 15243 9061 15255 9095
rect 15197 9055 15255 9061
rect 15378 9052 15384 9104
rect 15436 9052 15442 9104
rect 18138 9092 18144 9104
rect 16132 9064 18144 9092
rect 14458 8984 14464 9036
rect 14516 8984 14522 9036
rect 14734 8984 14740 9036
rect 14792 8984 14798 9036
rect 14829 9027 14887 9033
rect 14829 8993 14841 9027
rect 14875 8993 14887 9027
rect 14829 8987 14887 8993
rect 14844 8956 14872 8987
rect 14918 8984 14924 9036
rect 14976 8984 14982 9036
rect 15010 8984 15016 9036
rect 15068 9024 15074 9036
rect 16132 9033 16160 9064
rect 16117 9027 16175 9033
rect 16117 9024 16129 9027
rect 15068 8996 16129 9024
rect 15068 8984 15074 8996
rect 16117 8993 16129 8996
rect 16163 8993 16175 9027
rect 16117 8987 16175 8993
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 8993 16359 9027
rect 16301 8987 16359 8993
rect 15378 8956 15384 8968
rect 14384 8928 14688 8956
rect 14844 8928 15384 8956
rect 14553 8891 14611 8897
rect 14553 8888 14565 8891
rect 13740 8860 14565 8888
rect 11149 8823 11207 8829
rect 11149 8789 11161 8823
rect 11195 8789 11207 8823
rect 11149 8783 11207 8789
rect 11238 8780 11244 8832
rect 11296 8820 11302 8832
rect 11992 8829 12020 8860
rect 14553 8857 14565 8860
rect 14599 8857 14611 8891
rect 14553 8851 14611 8857
rect 11977 8823 12035 8829
rect 11977 8820 11989 8823
rect 11296 8792 11989 8820
rect 11296 8780 11302 8792
rect 11977 8789 11989 8792
rect 12023 8789 12035 8823
rect 11977 8783 12035 8789
rect 12434 8780 12440 8832
rect 12492 8780 12498 8832
rect 13446 8780 13452 8832
rect 13504 8780 13510 8832
rect 13906 8780 13912 8832
rect 13964 8780 13970 8832
rect 14090 8780 14096 8832
rect 14148 8780 14154 8832
rect 14660 8820 14688 8928
rect 15378 8916 15384 8928
rect 15436 8916 15442 8968
rect 15102 8848 15108 8900
rect 15160 8888 15166 8900
rect 15470 8888 15476 8900
rect 15160 8860 15476 8888
rect 15160 8848 15166 8860
rect 15470 8848 15476 8860
rect 15528 8848 15534 8900
rect 15194 8820 15200 8832
rect 14660 8792 15200 8820
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 15286 8780 15292 8832
rect 15344 8820 15350 8832
rect 15565 8823 15623 8829
rect 15565 8820 15577 8823
rect 15344 8792 15577 8820
rect 15344 8780 15350 8792
rect 15565 8789 15577 8792
rect 15611 8789 15623 8823
rect 16316 8820 16344 8987
rect 17586 8984 17592 9036
rect 17644 9033 17650 9036
rect 17880 9033 17908 9064
rect 18138 9052 18144 9064
rect 18196 9052 18202 9104
rect 18230 9052 18236 9104
rect 18288 9052 18294 9104
rect 18340 9092 18368 9132
rect 18443 9129 18455 9163
rect 18489 9160 18501 9163
rect 18782 9160 18788 9172
rect 18489 9132 18788 9160
rect 18489 9129 18501 9132
rect 18443 9123 18501 9129
rect 18782 9120 18788 9132
rect 18840 9120 18846 9172
rect 20162 9120 20168 9172
rect 20220 9120 20226 9172
rect 22554 9120 22560 9172
rect 22612 9160 22618 9172
rect 22741 9163 22799 9169
rect 22741 9160 22753 9163
rect 22612 9132 22753 9160
rect 22612 9120 22618 9132
rect 22741 9129 22753 9132
rect 22787 9129 22799 9163
rect 22741 9123 22799 9129
rect 20070 9092 20076 9104
rect 18340 9064 20076 9092
rect 20070 9052 20076 9064
rect 20128 9052 20134 9104
rect 20349 9095 20407 9101
rect 20349 9061 20361 9095
rect 20395 9092 20407 9095
rect 20438 9092 20444 9104
rect 20395 9064 20444 9092
rect 20395 9061 20407 9064
rect 20349 9055 20407 9061
rect 20438 9052 20444 9064
rect 20496 9052 20502 9104
rect 20530 9052 20536 9104
rect 20588 9092 20594 9104
rect 20901 9095 20959 9101
rect 20901 9092 20913 9095
rect 20588 9064 20913 9092
rect 20588 9052 20594 9064
rect 20901 9061 20913 9064
rect 20947 9092 20959 9095
rect 20947 9064 21128 9092
rect 20947 9061 20959 9064
rect 20901 9055 20959 9061
rect 17644 8987 17656 9033
rect 17865 9027 17923 9033
rect 17865 8993 17877 9027
rect 17911 8993 17923 9027
rect 18949 9027 19007 9033
rect 18949 9024 18961 9027
rect 17865 8987 17923 8993
rect 18616 8996 18961 9024
rect 17644 8984 17650 8987
rect 16390 8848 16396 8900
rect 16448 8888 16454 8900
rect 18616 8897 18644 8996
rect 18949 8993 18961 8996
rect 18995 8993 19007 9027
rect 18949 8987 19007 8993
rect 19242 8984 19248 9036
rect 19300 9024 19306 9036
rect 20162 9024 20168 9036
rect 19300 8996 20168 9024
rect 19300 8984 19306 8996
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 20254 8984 20260 9036
rect 20312 9024 20318 9036
rect 20622 9024 20628 9036
rect 20312 8996 20628 9024
rect 20312 8984 20318 8996
rect 20622 8984 20628 8996
rect 20680 9024 20686 9036
rect 20717 9027 20775 9033
rect 20717 9024 20729 9027
rect 20680 8996 20729 9024
rect 20680 8984 20686 8996
rect 20717 8993 20729 8996
rect 20763 8993 20775 9027
rect 21100 9024 21128 9064
rect 21266 9052 21272 9104
rect 21324 9092 21330 9104
rect 21606 9095 21664 9101
rect 21606 9092 21618 9095
rect 21324 9064 21618 9092
rect 21324 9052 21330 9064
rect 21606 9061 21618 9064
rect 21652 9061 21664 9095
rect 21606 9055 21664 9061
rect 22738 9024 22744 9036
rect 21100 8996 22744 9024
rect 20717 8987 20775 8993
rect 22738 8984 22744 8996
rect 22796 8984 22802 9036
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8925 18751 8959
rect 21085 8959 21143 8965
rect 21085 8956 21097 8959
rect 18693 8919 18751 8925
rect 19720 8928 21097 8956
rect 16485 8891 16543 8897
rect 16485 8888 16497 8891
rect 16448 8860 16497 8888
rect 16448 8848 16454 8860
rect 16485 8857 16497 8860
rect 16531 8857 16543 8891
rect 16485 8851 16543 8857
rect 18601 8891 18659 8897
rect 18601 8857 18613 8891
rect 18647 8857 18659 8891
rect 18601 8851 18659 8857
rect 18322 8820 18328 8832
rect 16316 8792 18328 8820
rect 15565 8783 15623 8789
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 18414 8780 18420 8832
rect 18472 8780 18478 8832
rect 18708 8820 18736 8919
rect 18874 8820 18880 8832
rect 18708 8792 18880 8820
rect 18874 8780 18880 8792
rect 18932 8820 18938 8832
rect 19720 8820 19748 8928
rect 21085 8925 21097 8928
rect 21131 8956 21143 8959
rect 21174 8956 21180 8968
rect 21131 8928 21180 8956
rect 21131 8925 21143 8928
rect 21085 8919 21143 8925
rect 21174 8916 21180 8928
rect 21232 8956 21238 8968
rect 21358 8956 21364 8968
rect 21232 8928 21364 8956
rect 21232 8916 21238 8928
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 19794 8848 19800 8900
rect 19852 8888 19858 8900
rect 20073 8891 20131 8897
rect 20073 8888 20085 8891
rect 19852 8860 20085 8888
rect 19852 8848 19858 8860
rect 20073 8857 20085 8860
rect 20119 8888 20131 8891
rect 20119 8860 21128 8888
rect 20119 8857 20131 8860
rect 20073 8851 20131 8857
rect 18932 8792 19748 8820
rect 18932 8780 18938 8792
rect 20162 8780 20168 8832
rect 20220 8820 20226 8832
rect 20349 8823 20407 8829
rect 20349 8820 20361 8823
rect 20220 8792 20361 8820
rect 20220 8780 20226 8792
rect 20349 8789 20361 8792
rect 20395 8820 20407 8823
rect 20714 8820 20720 8832
rect 20395 8792 20720 8820
rect 20395 8789 20407 8792
rect 20349 8783 20407 8789
rect 20714 8780 20720 8792
rect 20772 8820 20778 8832
rect 20990 8820 20996 8832
rect 20772 8792 20996 8820
rect 20772 8780 20778 8792
rect 20990 8780 20996 8792
rect 21048 8780 21054 8832
rect 21100 8820 21128 8860
rect 21542 8820 21548 8832
rect 21100 8792 21548 8820
rect 21542 8780 21548 8792
rect 21600 8780 21606 8832
rect 552 8730 23368 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 23368 8730
rect 552 8656 23368 8678
rect 7098 8576 7104 8628
rect 7156 8616 7162 8628
rect 7653 8619 7711 8625
rect 7653 8616 7665 8619
rect 7156 8588 7665 8616
rect 7156 8576 7162 8588
rect 7653 8585 7665 8588
rect 7699 8585 7711 8619
rect 7653 8579 7711 8585
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7892 8588 8033 8616
rect 7892 8576 7898 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 8386 8616 8392 8628
rect 8251 8588 8392 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 9953 8619 10011 8625
rect 9953 8616 9965 8619
rect 9824 8588 9965 8616
rect 9824 8576 9830 8588
rect 9953 8585 9965 8588
rect 9999 8585 10011 8619
rect 9953 8579 10011 8585
rect 10318 8576 10324 8628
rect 10376 8576 10382 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 12434 8616 12440 8628
rect 11195 8588 12440 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 12802 8576 12808 8628
rect 12860 8576 12866 8628
rect 13173 8619 13231 8625
rect 13173 8585 13185 8619
rect 13219 8616 13231 8619
rect 13633 8619 13691 8625
rect 13633 8616 13645 8619
rect 13219 8588 13645 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 13633 8585 13645 8588
rect 13679 8585 13691 8619
rect 15010 8616 15016 8628
rect 13633 8579 13691 8585
rect 13832 8588 15016 8616
rect 4890 8508 4896 8560
rect 4948 8548 4954 8560
rect 8294 8548 8300 8560
rect 4948 8520 8300 8548
rect 4948 8508 4954 8520
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 10137 8551 10195 8557
rect 10137 8517 10149 8551
rect 10183 8548 10195 8551
rect 11054 8548 11060 8560
rect 10183 8520 11060 8548
rect 10183 8517 10195 8520
rect 10137 8511 10195 8517
rect 11054 8508 11060 8520
rect 11112 8508 11118 8560
rect 11333 8551 11391 8557
rect 11333 8517 11345 8551
rect 11379 8517 11391 8551
rect 11333 8511 11391 8517
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8480 10839 8483
rect 11238 8480 11244 8492
rect 10827 8452 11244 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11348 8480 11376 8511
rect 11348 8452 11560 8480
rect 5626 8372 5632 8424
rect 5684 8412 5690 8424
rect 5905 8415 5963 8421
rect 5905 8412 5917 8415
rect 5684 8384 5917 8412
rect 5684 8372 5690 8384
rect 5905 8381 5917 8384
rect 5951 8381 5963 8415
rect 5905 8375 5963 8381
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8412 7619 8415
rect 7650 8412 7656 8424
rect 7607 8384 7656 8412
rect 7607 8381 7619 8384
rect 7561 8375 7619 8381
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 8478 8412 8484 8424
rect 7791 8384 8484 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 5721 8347 5779 8353
rect 5721 8313 5733 8347
rect 5767 8313 5779 8347
rect 5721 8307 5779 8313
rect 6089 8347 6147 8353
rect 6089 8313 6101 8347
rect 6135 8344 6147 8347
rect 7466 8344 7472 8356
rect 6135 8316 7472 8344
rect 6135 8313 6147 8316
rect 6089 8307 6147 8313
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 5736 8276 5764 8307
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 5994 8276 6000 8288
rect 4764 8248 6000 8276
rect 4764 8236 4770 8248
rect 5994 8236 6000 8248
rect 6052 8276 6058 8288
rect 6914 8276 6920 8288
rect 6052 8248 6920 8276
rect 6052 8236 6058 8248
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 7668 8276 7696 8372
rect 7760 8344 7788 8375
rect 8478 8372 8484 8384
rect 8536 8372 8542 8424
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 8662 8412 8668 8424
rect 8619 8384 8668 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 11330 8372 11336 8424
rect 11388 8412 11394 8424
rect 11425 8415 11483 8421
rect 11425 8412 11437 8415
rect 11388 8384 11437 8412
rect 11388 8372 11394 8384
rect 11425 8381 11437 8384
rect 11471 8381 11483 8415
rect 11532 8412 11560 8452
rect 11681 8415 11739 8421
rect 11681 8412 11693 8415
rect 11532 8384 11693 8412
rect 11425 8375 11483 8381
rect 11681 8381 11693 8384
rect 11727 8381 11739 8415
rect 11681 8375 11739 8381
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 7837 8347 7895 8353
rect 7837 8344 7849 8347
rect 7760 8316 7849 8344
rect 7837 8313 7849 8316
rect 7883 8313 7895 8347
rect 7837 8307 7895 8313
rect 8840 8347 8898 8353
rect 8840 8313 8852 8347
rect 8886 8344 8898 8347
rect 9306 8344 9312 8356
rect 8886 8316 9312 8344
rect 8886 8313 8898 8316
rect 8840 8307 8898 8313
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 10321 8347 10379 8353
rect 10321 8344 10333 8347
rect 10192 8316 10333 8344
rect 10192 8304 10198 8316
rect 10321 8313 10333 8316
rect 10367 8344 10379 8347
rect 11149 8347 11207 8353
rect 11149 8344 11161 8347
rect 10367 8316 11161 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 11149 8313 11161 8316
rect 11195 8344 11207 8347
rect 12986 8344 12992 8356
rect 11195 8316 12992 8344
rect 11195 8313 11207 8316
rect 11149 8307 11207 8313
rect 12986 8304 12992 8316
rect 13044 8304 13050 8356
rect 13205 8347 13263 8353
rect 13205 8313 13217 8347
rect 13251 8344 13263 8347
rect 13446 8344 13452 8356
rect 13251 8316 13452 8344
rect 13251 8313 13263 8316
rect 13205 8307 13263 8313
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 13556 8344 13584 8375
rect 13722 8372 13728 8424
rect 13780 8372 13786 8424
rect 13832 8421 13860 8588
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15378 8616 15384 8628
rect 15335 8588 15384 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 16390 8576 16396 8628
rect 16448 8616 16454 8628
rect 16448 8588 16804 8616
rect 16448 8576 16454 8588
rect 13817 8415 13875 8421
rect 13817 8381 13829 8415
rect 13863 8381 13875 8415
rect 13817 8375 13875 8381
rect 13906 8372 13912 8424
rect 13964 8412 13970 8424
rect 14073 8415 14131 8421
rect 14073 8412 14085 8415
rect 13964 8384 14085 8412
rect 13964 8372 13970 8384
rect 14073 8381 14085 8384
rect 14119 8381 14131 8415
rect 14073 8375 14131 8381
rect 15010 8372 15016 8424
rect 15068 8412 15074 8424
rect 16669 8415 16727 8421
rect 16669 8412 16681 8415
rect 15068 8384 16681 8412
rect 15068 8372 15074 8384
rect 16669 8381 16681 8384
rect 16715 8381 16727 8415
rect 16776 8412 16804 8588
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 16908 8588 17417 8616
rect 16908 8576 16914 8588
rect 17405 8585 17417 8588
rect 17451 8585 17463 8619
rect 17405 8579 17463 8585
rect 17586 8576 17592 8628
rect 17644 8576 17650 8628
rect 18322 8576 18328 8628
rect 18380 8616 18386 8628
rect 19978 8616 19984 8628
rect 18380 8588 19984 8616
rect 18380 8576 18386 8588
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 20438 8576 20444 8628
rect 20496 8576 20502 8628
rect 21729 8619 21787 8625
rect 21729 8616 21741 8619
rect 20824 8588 21741 8616
rect 20824 8560 20852 8588
rect 21729 8585 21741 8588
rect 21775 8585 21787 8619
rect 21729 8579 21787 8585
rect 22189 8619 22247 8625
rect 22189 8585 22201 8619
rect 22235 8616 22247 8619
rect 22370 8616 22376 8628
rect 22235 8588 22376 8616
rect 22235 8585 22247 8588
rect 22189 8579 22247 8585
rect 22370 8576 22376 8588
rect 22428 8576 22434 8628
rect 22465 8619 22523 8625
rect 22465 8585 22477 8619
rect 22511 8616 22523 8619
rect 22554 8616 22560 8628
rect 22511 8588 22560 8616
rect 22511 8585 22523 8588
rect 22465 8579 22523 8585
rect 22554 8576 22560 8588
rect 22612 8576 22618 8628
rect 19886 8508 19892 8560
rect 19944 8548 19950 8560
rect 20257 8551 20315 8557
rect 20257 8548 20269 8551
rect 19944 8520 20269 8548
rect 19944 8508 19950 8520
rect 20257 8517 20269 8520
rect 20303 8517 20315 8551
rect 20806 8548 20812 8560
rect 20257 8511 20315 8517
rect 20640 8520 20812 8548
rect 18874 8440 18880 8492
rect 18932 8440 18938 8492
rect 19150 8421 19156 8424
rect 16945 8415 17003 8421
rect 16945 8412 16957 8415
rect 16776 8384 16957 8412
rect 16669 8375 16727 8381
rect 16945 8381 16957 8384
rect 16991 8381 17003 8415
rect 16945 8375 17003 8381
rect 17129 8415 17187 8421
rect 17129 8381 17141 8415
rect 17175 8412 17187 8415
rect 19144 8412 19156 8421
rect 17175 8384 17356 8412
rect 19111 8384 19156 8412
rect 17175 8381 17187 8384
rect 17129 8375 17187 8381
rect 14918 8344 14924 8356
rect 13556 8316 14924 8344
rect 14918 8304 14924 8316
rect 14976 8304 14982 8356
rect 15470 8304 15476 8356
rect 15528 8344 15534 8356
rect 16402 8347 16460 8353
rect 16402 8344 16414 8347
rect 15528 8316 16414 8344
rect 15528 8304 15534 8316
rect 16402 8313 16414 8316
rect 16448 8313 16460 8347
rect 16402 8307 16460 8313
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 16761 8347 16819 8353
rect 16761 8344 16773 8347
rect 16632 8316 16773 8344
rect 16632 8304 16638 8316
rect 16761 8313 16773 8316
rect 16807 8313 16819 8347
rect 17218 8344 17224 8356
rect 16761 8307 16819 8313
rect 16868 8316 17224 8344
rect 8037 8279 8095 8285
rect 8037 8276 8049 8279
rect 7668 8248 8049 8276
rect 8037 8245 8049 8248
rect 8083 8245 8095 8279
rect 8037 8239 8095 8245
rect 13354 8236 13360 8288
rect 13412 8236 13418 8288
rect 14274 8236 14280 8288
rect 14332 8276 14338 8288
rect 14734 8276 14740 8288
rect 14332 8248 14740 8276
rect 14332 8236 14338 8248
rect 14734 8236 14740 8248
rect 14792 8276 14798 8288
rect 15197 8279 15255 8285
rect 15197 8276 15209 8279
rect 14792 8248 15209 8276
rect 14792 8236 14798 8248
rect 15197 8245 15209 8248
rect 15243 8245 15255 8279
rect 15197 8239 15255 8245
rect 15378 8236 15384 8288
rect 15436 8276 15442 8288
rect 16868 8276 16896 8316
rect 17218 8304 17224 8316
rect 17276 8304 17282 8356
rect 17328 8344 17356 8384
rect 19144 8375 19156 8384
rect 19150 8372 19156 8375
rect 19208 8372 19214 8424
rect 20640 8421 20668 8520
rect 20806 8508 20812 8520
rect 20864 8508 20870 8560
rect 21910 8548 21916 8560
rect 21284 8520 21916 8548
rect 20625 8415 20683 8421
rect 20625 8381 20637 8415
rect 20671 8381 20683 8415
rect 20885 8415 20943 8421
rect 20885 8412 20897 8415
rect 20625 8375 20683 8381
rect 20824 8384 20897 8412
rect 17421 8347 17479 8353
rect 17421 8344 17433 8347
rect 17328 8316 17433 8344
rect 17421 8313 17433 8316
rect 17467 8313 17479 8347
rect 17421 8307 17479 8313
rect 20714 8304 20720 8356
rect 20772 8344 20778 8356
rect 20824 8344 20852 8384
rect 20885 8381 20897 8384
rect 20931 8381 20943 8415
rect 20885 8375 20943 8381
rect 20990 8372 20996 8424
rect 21048 8372 21054 8424
rect 21174 8372 21180 8424
rect 21232 8372 21238 8424
rect 21284 8421 21312 8520
rect 21910 8508 21916 8520
rect 21968 8548 21974 8560
rect 22281 8551 22339 8557
rect 22281 8548 22293 8551
rect 21968 8520 22293 8548
rect 21968 8508 21974 8520
rect 22281 8517 22293 8520
rect 22327 8517 22339 8551
rect 22281 8511 22339 8517
rect 22738 8508 22744 8560
rect 22796 8508 22802 8560
rect 21450 8440 21456 8492
rect 21508 8480 21514 8492
rect 21508 8452 21579 8480
rect 21508 8440 21514 8452
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8381 21327 8415
rect 21269 8375 21327 8381
rect 21361 8415 21419 8421
rect 21361 8381 21373 8415
rect 21407 8409 21419 8415
rect 21468 8409 21496 8440
rect 21407 8381 21496 8409
rect 21551 8412 21579 8452
rect 21634 8440 21640 8492
rect 21692 8440 21698 8492
rect 21818 8440 21824 8492
rect 21876 8440 21882 8492
rect 22002 8412 22008 8424
rect 21551 8384 22008 8412
rect 21361 8375 21419 8381
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 22922 8372 22928 8424
rect 22980 8372 22986 8424
rect 20772 8316 20852 8344
rect 20772 8304 20778 8316
rect 21542 8304 21548 8356
rect 21600 8344 21606 8356
rect 21729 8347 21787 8353
rect 21729 8344 21741 8347
rect 21600 8316 21741 8344
rect 21600 8304 21606 8316
rect 21729 8313 21741 8316
rect 21775 8313 21787 8347
rect 21729 8307 21787 8313
rect 22186 8304 22192 8356
rect 22244 8344 22250 8356
rect 22433 8347 22491 8353
rect 22433 8344 22445 8347
rect 22244 8316 22445 8344
rect 22244 8304 22250 8316
rect 22433 8313 22445 8316
rect 22479 8313 22491 8347
rect 22433 8307 22491 8313
rect 22646 8304 22652 8356
rect 22704 8304 22710 8356
rect 15436 8248 16896 8276
rect 20809 8279 20867 8285
rect 15436 8236 15442 8248
rect 20809 8245 20821 8279
rect 20855 8276 20867 8279
rect 20898 8276 20904 8288
rect 20855 8248 20904 8276
rect 20855 8245 20867 8248
rect 20809 8239 20867 8245
rect 20898 8236 20904 8248
rect 20956 8276 20962 8288
rect 21450 8276 21456 8288
rect 20956 8248 21456 8276
rect 20956 8236 20962 8248
rect 21450 8236 21456 8248
rect 21508 8236 21514 8288
rect 552 8186 23368 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 23368 8186
rect 552 8112 23368 8134
rect 5077 8075 5135 8081
rect 5077 8041 5089 8075
rect 5123 8072 5135 8075
rect 5902 8072 5908 8084
rect 5123 8044 5908 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 7834 8032 7840 8084
rect 7892 8032 7898 8084
rect 8202 8032 8208 8084
rect 8260 8072 8266 8084
rect 8260 8044 9168 8072
rect 8260 8032 8266 8044
rect 4430 7964 4436 8016
rect 4488 8004 4494 8016
rect 4709 8007 4767 8013
rect 4709 8004 4721 8007
rect 4488 7976 4721 8004
rect 4488 7964 4494 7976
rect 4709 7973 4721 7976
rect 4755 7973 4767 8007
rect 4709 7967 4767 7973
rect 4925 8007 4983 8013
rect 4925 7973 4937 8007
rect 4971 8004 4983 8007
rect 6457 8007 6515 8013
rect 6457 8004 6469 8007
rect 4971 7976 6469 8004
rect 4971 7973 4983 7976
rect 4925 7967 4983 7973
rect 6457 7973 6469 7976
rect 6503 7973 6515 8007
rect 6457 7967 6515 7973
rect 8938 7964 8944 8016
rect 8996 8013 9002 8016
rect 8996 8004 9008 8013
rect 9140 8004 9168 8044
rect 9306 8032 9312 8084
rect 9364 8032 9370 8084
rect 10318 8032 10324 8084
rect 10376 8032 10382 8084
rect 11606 8072 11612 8084
rect 10520 8044 11612 8072
rect 9493 8007 9551 8013
rect 9493 8004 9505 8007
rect 8996 7976 9041 8004
rect 9140 7976 9505 8004
rect 8996 7967 9008 7976
rect 9493 7973 9505 7976
rect 9539 8004 9551 8007
rect 9953 8007 10011 8013
rect 9953 8004 9965 8007
rect 9539 7976 9965 8004
rect 9539 7973 9551 7976
rect 9493 7967 9551 7973
rect 9953 7973 9965 7976
rect 9999 7973 10011 8007
rect 9953 7967 10011 7973
rect 8996 7964 9002 7967
rect 10134 7964 10140 8016
rect 10192 7964 10198 8016
rect 4522 7896 4528 7948
rect 4580 7936 4586 7948
rect 5997 7939 6055 7945
rect 5997 7936 6009 7939
rect 4580 7908 6009 7936
rect 4580 7896 4586 7908
rect 5997 7905 6009 7908
rect 6043 7936 6055 7939
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 6043 7908 6653 7936
rect 6043 7905 6055 7908
rect 5997 7899 6055 7905
rect 6641 7905 6653 7908
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 5074 7828 5080 7880
rect 5132 7868 5138 7880
rect 5132 7840 5396 7868
rect 5132 7828 5138 7840
rect 4982 7800 4988 7812
rect 4908 7772 4988 7800
rect 4908 7741 4936 7772
rect 4982 7760 4988 7772
rect 5040 7800 5046 7812
rect 5258 7800 5264 7812
rect 5040 7772 5264 7800
rect 5040 7760 5046 7772
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 4893 7735 4951 7741
rect 4893 7701 4905 7735
rect 4939 7701 4951 7735
rect 4893 7695 4951 7701
rect 5166 7692 5172 7744
rect 5224 7692 5230 7744
rect 5368 7732 5396 7840
rect 5626 7828 5632 7880
rect 5684 7828 5690 7880
rect 6086 7828 6092 7880
rect 6144 7828 6150 7880
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7837 6239 7871
rect 6181 7831 6239 7837
rect 5644 7800 5672 7828
rect 5644 7772 5948 7800
rect 5813 7735 5871 7741
rect 5813 7732 5825 7735
rect 5368 7704 5825 7732
rect 5813 7701 5825 7704
rect 5859 7701 5871 7735
rect 5920 7732 5948 7772
rect 6196 7732 6224 7831
rect 6270 7828 6276 7880
rect 6328 7828 6334 7880
rect 6656 7800 6684 7899
rect 6822 7896 6828 7948
rect 6880 7896 6886 7948
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7098 7936 7104 7948
rect 6972 7908 7104 7936
rect 6972 7896 6978 7908
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 8662 7896 8668 7948
rect 8720 7936 8726 7948
rect 10520 7945 10548 8044
rect 11606 8032 11612 8044
rect 11664 8072 11670 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 11664 8044 12357 8072
rect 11664 8032 11670 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 12345 8035 12403 8041
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 14458 8072 14464 8084
rect 13872 8044 14464 8072
rect 13872 8032 13878 8044
rect 14458 8032 14464 8044
rect 14516 8072 14522 8084
rect 14737 8075 14795 8081
rect 14737 8072 14749 8075
rect 14516 8044 14749 8072
rect 14516 8032 14522 8044
rect 14737 8041 14749 8044
rect 14783 8041 14795 8075
rect 14737 8035 14795 8041
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 15289 8075 15347 8081
rect 15289 8072 15301 8075
rect 15252 8044 15301 8072
rect 15252 8032 15258 8044
rect 15289 8041 15301 8044
rect 15335 8072 15347 8075
rect 15378 8072 15384 8084
rect 15335 8044 15384 8072
rect 15335 8041 15347 8044
rect 15289 8035 15347 8041
rect 15378 8032 15384 8044
rect 15436 8032 15442 8084
rect 15470 8032 15476 8084
rect 15528 8032 15534 8084
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 19245 8075 19303 8081
rect 19245 8072 19257 8075
rect 18472 8044 19257 8072
rect 18472 8032 18478 8044
rect 19245 8041 19257 8044
rect 19291 8041 19303 8075
rect 19245 8035 19303 8041
rect 19702 8032 19708 8084
rect 19760 8032 19766 8084
rect 20622 8072 20628 8084
rect 20088 8044 20628 8072
rect 10689 8007 10747 8013
rect 10689 7973 10701 8007
rect 10735 8004 10747 8007
rect 10870 8004 10876 8016
rect 10735 7976 10876 8004
rect 10735 7973 10747 7976
rect 10689 7967 10747 7973
rect 10870 7964 10876 7976
rect 10928 7964 10934 8016
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 11210 8007 11268 8013
rect 11210 8004 11222 8007
rect 11112 7976 11222 8004
rect 11112 7964 11118 7976
rect 11210 7973 11222 7976
rect 11256 7973 11268 8007
rect 11210 7967 11268 7973
rect 11330 7964 11336 8016
rect 11388 8004 11394 8016
rect 13265 8007 13323 8013
rect 13265 8004 13277 8007
rect 11388 7976 13277 8004
rect 11388 7964 11394 7976
rect 13265 7973 13277 7976
rect 13311 7973 13323 8007
rect 13265 7967 13323 7973
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 8720 7908 9229 7936
rect 8720 7896 8726 7908
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 10505 7939 10563 7945
rect 10505 7905 10517 7939
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 10778 7896 10784 7948
rect 10836 7896 10842 7948
rect 13078 7896 13084 7948
rect 13136 7896 13142 7948
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7868 9919 7871
rect 10796 7868 10824 7896
rect 9907 7840 10824 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 10962 7828 10968 7880
rect 11020 7828 11026 7880
rect 13280 7868 13308 7967
rect 13354 7964 13360 8016
rect 13412 8004 13418 8016
rect 13602 8007 13660 8013
rect 13602 8004 13614 8007
rect 13412 7976 13614 8004
rect 13412 7964 13418 7976
rect 13602 7973 13614 7976
rect 13648 7973 13660 8007
rect 13602 7967 13660 7973
rect 19610 7964 19616 8016
rect 19668 7964 19674 8016
rect 19886 7964 19892 8016
rect 19944 7964 19950 8016
rect 20088 8013 20116 8044
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 21910 8072 21916 8084
rect 20808 8044 21916 8072
rect 20073 8007 20131 8013
rect 20073 7973 20085 8007
rect 20119 7973 20131 8007
rect 20073 7967 20131 7973
rect 20714 7964 20720 8016
rect 20772 8004 20778 8016
rect 20808 8004 20836 8044
rect 21910 8032 21916 8044
rect 21968 8032 21974 8084
rect 22002 8032 22008 8084
rect 22060 8072 22066 8084
rect 22649 8075 22707 8081
rect 22649 8072 22661 8075
rect 22060 8044 22661 8072
rect 22060 8032 22066 8044
rect 22649 8041 22661 8044
rect 22695 8041 22707 8075
rect 22649 8035 22707 8041
rect 20772 7973 20836 8004
rect 20772 7964 20775 7973
rect 14921 7939 14979 7945
rect 14921 7905 14933 7939
rect 14967 7936 14979 7939
rect 15102 7936 15108 7948
rect 14967 7908 15108 7936
rect 14967 7905 14979 7908
rect 14921 7899 14979 7905
rect 15102 7896 15108 7908
rect 15160 7896 15166 7948
rect 19429 7939 19487 7945
rect 19429 7905 19441 7939
rect 19475 7936 19487 7939
rect 19794 7936 19800 7948
rect 19475 7908 19800 7936
rect 19475 7905 19487 7908
rect 19429 7899 19487 7905
rect 19794 7896 19800 7908
rect 19852 7896 19858 7948
rect 20763 7939 20775 7964
rect 20809 7942 20836 7973
rect 20898 7964 20904 8016
rect 20956 8004 20962 8016
rect 20993 8007 21051 8013
rect 20993 8004 21005 8007
rect 20956 7976 21005 8004
rect 20956 7964 20962 7976
rect 20993 7973 21005 7976
rect 21039 7973 21051 8007
rect 20993 7967 21051 7973
rect 21536 8007 21594 8013
rect 21536 7973 21548 8007
rect 21582 8004 21594 8007
rect 21634 8004 21640 8016
rect 21582 7976 21640 8004
rect 21582 7973 21594 7976
rect 21536 7967 21594 7973
rect 21634 7964 21640 7976
rect 21692 7964 21698 8016
rect 20809 7939 20821 7942
rect 20763 7933 20821 7939
rect 21358 7896 21364 7948
rect 21416 7896 21422 7948
rect 13357 7871 13415 7877
rect 13357 7868 13369 7871
rect 13280 7840 13369 7868
rect 13357 7837 13369 7840
rect 13403 7837 13415 7871
rect 13357 7831 13415 7837
rect 21269 7871 21327 7877
rect 21269 7837 21281 7871
rect 21315 7868 21327 7871
rect 21376 7868 21404 7896
rect 21315 7840 21404 7868
rect 21315 7837 21327 7840
rect 21269 7831 21327 7837
rect 6914 7800 6920 7812
rect 6656 7772 6920 7800
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 6822 7732 6828 7744
rect 5920 7704 6828 7732
rect 5813 7695 5871 7701
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 9490 7692 9496 7744
rect 9548 7692 9554 7744
rect 15286 7692 15292 7744
rect 15344 7692 15350 7744
rect 20806 7692 20812 7744
rect 20864 7692 20870 7744
rect 552 7642 23368 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 23368 7642
rect 552 7568 23368 7590
rect 4430 7488 4436 7540
rect 4488 7488 4494 7540
rect 4982 7488 4988 7540
rect 5040 7488 5046 7540
rect 6270 7488 6276 7540
rect 6328 7528 6334 7540
rect 6641 7531 6699 7537
rect 6641 7528 6653 7531
rect 6328 7500 6653 7528
rect 6328 7488 6334 7500
rect 6641 7497 6653 7500
rect 6687 7497 6699 7531
rect 6641 7491 6699 7497
rect 7561 7531 7619 7537
rect 7561 7497 7573 7531
rect 7607 7528 7619 7531
rect 8202 7528 8208 7540
rect 7607 7500 8208 7528
rect 7607 7497 7619 7500
rect 7561 7491 7619 7497
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7392 4675 7395
rect 4663 7364 5396 7392
rect 4663 7361 4675 7364
rect 4617 7355 4675 7361
rect 5368 7336 5396 7364
rect 4246 7284 4252 7336
rect 4304 7284 4310 7336
rect 4522 7284 4528 7336
rect 4580 7284 4586 7336
rect 5258 7284 5264 7336
rect 5316 7284 5322 7336
rect 5350 7284 5356 7336
rect 5408 7324 5414 7336
rect 6656 7324 6684 7491
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 11609 7531 11667 7537
rect 11609 7528 11621 7531
rect 10928 7500 11621 7528
rect 10928 7488 10934 7500
rect 11609 7497 11621 7500
rect 11655 7497 11667 7531
rect 11609 7491 11667 7497
rect 14090 7488 14096 7540
rect 14148 7488 14154 7540
rect 21174 7488 21180 7540
rect 21232 7488 21238 7540
rect 6822 7420 6828 7472
rect 6880 7460 6886 7472
rect 7285 7463 7343 7469
rect 7285 7460 7297 7463
rect 6880 7432 7297 7460
rect 6880 7420 6886 7432
rect 7285 7429 7297 7432
rect 7331 7429 7343 7463
rect 7285 7423 7343 7429
rect 8662 7420 8668 7472
rect 8720 7420 8726 7472
rect 7009 7327 7067 7333
rect 7009 7324 7021 7327
rect 5408 7296 5672 7324
rect 6656 7296 7021 7324
rect 5408 7284 5414 7296
rect 4341 7259 4399 7265
rect 4341 7225 4353 7259
rect 4387 7256 4399 7259
rect 4706 7256 4712 7268
rect 4387 7228 4712 7256
rect 4387 7225 4399 7228
rect 4341 7219 4399 7225
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 4985 7259 5043 7265
rect 4985 7225 4997 7259
rect 5031 7256 5043 7259
rect 5074 7256 5080 7268
rect 5031 7228 5080 7256
rect 5031 7225 5043 7228
rect 4985 7219 5043 7225
rect 5074 7216 5080 7228
rect 5132 7216 5138 7268
rect 5506 7259 5564 7265
rect 5506 7256 5518 7259
rect 5184 7228 5518 7256
rect 5184 7197 5212 7228
rect 5506 7225 5518 7228
rect 5552 7225 5564 7259
rect 5644 7256 5672 7296
rect 7009 7293 7021 7296
rect 7055 7293 7067 7327
rect 7009 7287 7067 7293
rect 7098 7284 7104 7336
rect 7156 7284 7162 7336
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 8352 7296 8861 7324
rect 8352 7284 8358 7296
rect 8849 7293 8861 7296
rect 8895 7324 8907 7327
rect 10229 7327 10287 7333
rect 10229 7324 10241 7327
rect 8895 7296 10241 7324
rect 8895 7293 8907 7296
rect 8849 7287 8907 7293
rect 10229 7293 10241 7296
rect 10275 7324 10287 7327
rect 11054 7324 11060 7336
rect 10275 7296 11060 7324
rect 10275 7293 10287 7296
rect 10229 7287 10287 7293
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 14274 7284 14280 7336
rect 14332 7284 14338 7336
rect 14458 7284 14464 7336
rect 14516 7284 14522 7336
rect 14553 7327 14611 7333
rect 14553 7293 14565 7327
rect 14599 7324 14611 7327
rect 14918 7324 14924 7336
rect 14599 7296 14924 7324
rect 14599 7293 14611 7296
rect 14553 7287 14611 7293
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 20898 7284 20904 7336
rect 20956 7324 20962 7336
rect 21085 7327 21143 7333
rect 21085 7324 21097 7327
rect 20956 7296 21097 7324
rect 20956 7284 20962 7296
rect 21085 7293 21097 7296
rect 21131 7293 21143 7327
rect 21085 7287 21143 7293
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 21910 7324 21916 7336
rect 21315 7296 21916 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 21910 7284 21916 7296
rect 21968 7284 21974 7336
rect 6733 7259 6791 7265
rect 6733 7256 6745 7259
rect 5644 7228 6745 7256
rect 5506 7219 5564 7225
rect 6733 7225 6745 7228
rect 6779 7225 6791 7259
rect 6733 7219 6791 7225
rect 6914 7216 6920 7268
rect 6972 7216 6978 7268
rect 7466 7216 7472 7268
rect 7524 7265 7530 7268
rect 7524 7259 7587 7265
rect 7524 7225 7541 7259
rect 7575 7225 7587 7259
rect 7524 7219 7587 7225
rect 7524 7216 7530 7219
rect 7742 7216 7748 7268
rect 7800 7216 7806 7268
rect 10496 7259 10554 7265
rect 10496 7225 10508 7259
rect 10542 7225 10554 7259
rect 10496 7219 10554 7225
rect 5169 7191 5227 7197
rect 5169 7157 5181 7191
rect 5215 7157 5227 7191
rect 5169 7151 5227 7157
rect 7374 7148 7380 7200
rect 7432 7148 7438 7200
rect 10410 7148 10416 7200
rect 10468 7188 10474 7200
rect 10520 7188 10548 7219
rect 10468 7160 10548 7188
rect 10468 7148 10474 7160
rect 552 7098 23368 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 23368 7098
rect 552 7024 23368 7046
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 5626 6984 5632 6996
rect 4304 6956 5632 6984
rect 4304 6944 4310 6956
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7193 6987 7251 6993
rect 7193 6984 7205 6987
rect 6972 6956 7205 6984
rect 6972 6944 6978 6956
rect 7193 6953 7205 6956
rect 7239 6953 7251 6987
rect 7193 6947 7251 6953
rect 7469 6987 7527 6993
rect 7469 6953 7481 6987
rect 7515 6984 7527 6987
rect 7742 6984 7748 6996
rect 7515 6956 7748 6984
rect 7515 6953 7527 6956
rect 7469 6947 7527 6953
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 10410 6944 10416 6996
rect 10468 6944 10474 6996
rect 10594 6993 10600 6996
rect 10581 6987 10600 6993
rect 10581 6953 10593 6987
rect 10581 6947 10600 6953
rect 10594 6944 10600 6947
rect 10652 6944 10658 6996
rect 5166 6876 5172 6928
rect 5224 6916 5230 6928
rect 5362 6919 5420 6925
rect 5362 6916 5374 6919
rect 5224 6888 5374 6916
rect 5224 6876 5230 6888
rect 5362 6885 5374 6888
rect 5408 6885 5420 6919
rect 5362 6879 5420 6885
rect 6822 6876 6828 6928
rect 6880 6916 6886 6928
rect 6880 6888 7512 6916
rect 6880 6876 6886 6888
rect 5902 6808 5908 6860
rect 5960 6848 5966 6860
rect 6069 6851 6127 6857
rect 6069 6848 6081 6851
rect 5960 6820 6081 6848
rect 5960 6808 5966 6820
rect 6069 6817 6081 6820
rect 6115 6817 6127 6851
rect 6069 6811 6127 6817
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 7484 6857 7512 6888
rect 10134 6876 10140 6928
rect 10192 6916 10198 6928
rect 10781 6919 10839 6925
rect 10781 6916 10793 6919
rect 10192 6888 10793 6916
rect 10192 6876 10198 6888
rect 10781 6885 10793 6888
rect 10827 6885 10839 6919
rect 10781 6879 10839 6885
rect 7285 6851 7343 6857
rect 7285 6848 7297 6851
rect 7156 6820 7297 6848
rect 7156 6808 7162 6820
rect 7285 6817 7297 6820
rect 7331 6817 7343 6851
rect 7285 6811 7343 6817
rect 7469 6851 7527 6857
rect 7469 6817 7481 6851
rect 7515 6817 7527 6851
rect 7469 6811 7527 6817
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6780 5687 6783
rect 5810 6780 5816 6792
rect 5675 6752 5816 6780
rect 5675 6749 5687 6752
rect 5629 6743 5687 6749
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5644 6644 5672 6743
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 5316 6616 5672 6644
rect 5316 6604 5322 6616
rect 10226 6604 10232 6656
rect 10284 6644 10290 6656
rect 10597 6647 10655 6653
rect 10597 6644 10609 6647
rect 10284 6616 10609 6644
rect 10284 6604 10290 6616
rect 10597 6613 10609 6616
rect 10643 6613 10655 6647
rect 10597 6607 10655 6613
rect 552 6554 23368 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 23368 6554
rect 552 6480 23368 6502
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 4764 6412 5457 6440
rect 4764 6400 4770 6412
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 5868 6412 6868 6440
rect 5868 6400 5874 6412
rect 6840 6313 6868 6412
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6304 6883 6307
rect 8662 6304 8668 6316
rect 6871 6276 8668 6304
rect 6871 6273 6883 6276
rect 6825 6267 6883 6273
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 6580 6171 6638 6177
rect 6580 6137 6592 6171
rect 6626 6168 6638 6171
rect 7374 6168 7380 6180
rect 6626 6140 7380 6168
rect 6626 6137 6638 6140
rect 6580 6131 6638 6137
rect 7374 6128 7380 6140
rect 7432 6128 7438 6180
rect 552 6010 23368 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 23368 6010
rect 552 5936 23368 5958
rect 552 5466 23368 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 23368 5466
rect 552 5392 23368 5414
rect 552 4922 23368 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 23368 4922
rect 552 4848 23368 4870
rect 552 4378 23368 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 23368 4378
rect 552 4304 23368 4326
rect 22833 4267 22891 4273
rect 22833 4233 22845 4267
rect 22879 4264 22891 4267
rect 22922 4264 22928 4276
rect 22879 4236 22928 4264
rect 22879 4233 22891 4236
rect 22833 4227 22891 4233
rect 22922 4224 22928 4236
rect 22980 4224 22986 4276
rect 23014 4020 23020 4072
rect 23072 4020 23078 4072
rect 552 3834 23368 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 23368 3834
rect 552 3760 23368 3782
rect 552 3290 23368 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 23368 3290
rect 552 3216 23368 3238
rect 552 2746 23368 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 23368 2746
rect 552 2672 23368 2694
rect 552 2202 23368 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 23368 2202
rect 552 2128 23368 2150
rect 552 1658 23368 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 23368 1658
rect 552 1584 23368 1606
rect 552 1114 23368 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 23368 1114
rect 552 1040 23368 1062
rect 552 570 23368 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 23368 570
rect 552 496 23368 518
<< via1 >>
rect 4322 23366 4374 23418
rect 4386 23366 4438 23418
rect 4450 23366 4502 23418
rect 4514 23366 4566 23418
rect 4578 23366 4630 23418
rect 7564 23264 7616 23316
rect 7656 23264 7708 23316
rect 19708 23264 19760 23316
rect 1768 23171 1820 23180
rect 1768 23137 1777 23171
rect 1777 23137 1811 23171
rect 1811 23137 1820 23171
rect 1768 23128 1820 23137
rect 4712 23171 4764 23180
rect 4712 23137 4721 23171
rect 4721 23137 4755 23171
rect 4755 23137 4764 23171
rect 4712 23128 4764 23137
rect 6276 23171 6328 23180
rect 6276 23137 6285 23171
rect 6285 23137 6319 23171
rect 6319 23137 6328 23171
rect 6276 23128 6328 23137
rect 7380 23128 7432 23180
rect 10416 23239 10468 23248
rect 10416 23205 10425 23239
rect 10425 23205 10459 23239
rect 10459 23205 10468 23239
rect 10416 23196 10468 23205
rect 6920 23060 6972 23112
rect 7656 23060 7708 23112
rect 5448 22992 5500 23044
rect 6184 22992 6236 23044
rect 9220 23128 9272 23180
rect 11060 23171 11112 23180
rect 11060 23137 11069 23171
rect 11069 23137 11103 23171
rect 11103 23137 11112 23171
rect 11060 23128 11112 23137
rect 11244 23128 11296 23180
rect 9588 23060 9640 23112
rect 10968 23060 11020 23112
rect 11888 23128 11940 23180
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 14464 23196 14516 23248
rect 18144 23196 18196 23248
rect 18696 23196 18748 23248
rect 15108 23128 15160 23180
rect 16396 23128 16448 23180
rect 18420 23128 18472 23180
rect 19524 23239 19576 23248
rect 19524 23205 19533 23239
rect 19533 23205 19567 23239
rect 19567 23205 19576 23239
rect 19524 23196 19576 23205
rect 19892 23239 19944 23248
rect 19892 23205 19901 23239
rect 19901 23205 19935 23239
rect 19935 23205 19944 23239
rect 19892 23196 19944 23205
rect 20076 23196 20128 23248
rect 18788 23103 18840 23112
rect 18788 23069 18797 23103
rect 18797 23069 18831 23103
rect 18831 23069 18840 23103
rect 18788 23060 18840 23069
rect 19064 23128 19116 23180
rect 20996 23196 21048 23248
rect 19892 23060 19944 23112
rect 9404 22992 9456 23044
rect 16028 22992 16080 23044
rect 21088 23128 21140 23180
rect 21364 23171 21416 23180
rect 21364 23137 21373 23171
rect 21373 23137 21407 23171
rect 21407 23137 21416 23171
rect 21364 23128 21416 23137
rect 21456 23128 21508 23180
rect 20536 23060 20588 23112
rect 21916 23171 21968 23180
rect 21916 23137 21925 23171
rect 21925 23137 21959 23171
rect 21959 23137 21968 23171
rect 21916 23128 21968 23137
rect 22284 23128 22336 23180
rect 4896 22967 4948 22976
rect 4896 22933 4905 22967
rect 4905 22933 4939 22967
rect 4939 22933 4948 22967
rect 4896 22924 4948 22933
rect 5356 22924 5408 22976
rect 7748 22924 7800 22976
rect 13544 22924 13596 22976
rect 14280 22924 14332 22976
rect 17500 22924 17552 22976
rect 19984 22967 20036 22976
rect 19984 22933 19993 22967
rect 19993 22933 20027 22967
rect 20027 22933 20036 22967
rect 19984 22924 20036 22933
rect 20076 22924 20128 22976
rect 21364 22924 21416 22976
rect 21732 22924 21784 22976
rect 22560 22924 22612 22976
rect 3662 22822 3714 22874
rect 3726 22822 3778 22874
rect 3790 22822 3842 22874
rect 3854 22822 3906 22874
rect 3918 22822 3970 22874
rect 9772 22720 9824 22772
rect 10416 22720 10468 22772
rect 14004 22720 14056 22772
rect 14280 22763 14332 22772
rect 14280 22729 14289 22763
rect 14289 22729 14323 22763
rect 14323 22729 14332 22763
rect 14280 22720 14332 22729
rect 15200 22720 15252 22772
rect 5356 22652 5408 22704
rect 7380 22652 7432 22704
rect 9956 22652 10008 22704
rect 11060 22652 11112 22704
rect 4896 22584 4948 22636
rect 5632 22584 5684 22636
rect 4896 22491 4948 22500
rect 4896 22457 4905 22491
rect 4905 22457 4939 22491
rect 4939 22457 4948 22491
rect 4896 22448 4948 22457
rect 5448 22559 5500 22568
rect 5448 22525 5457 22559
rect 5457 22525 5491 22559
rect 5491 22525 5500 22559
rect 5448 22516 5500 22525
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 6368 22559 6420 22568
rect 6368 22525 6377 22559
rect 6377 22525 6411 22559
rect 6411 22525 6420 22559
rect 6368 22516 6420 22525
rect 7196 22559 7248 22568
rect 7196 22525 7205 22559
rect 7205 22525 7239 22559
rect 7239 22525 7248 22559
rect 7196 22516 7248 22525
rect 9220 22559 9272 22568
rect 9220 22525 9229 22559
rect 9229 22525 9263 22559
rect 9263 22525 9272 22559
rect 9220 22516 9272 22525
rect 6000 22448 6052 22500
rect 6184 22491 6236 22500
rect 6184 22457 6193 22491
rect 6193 22457 6227 22491
rect 6227 22457 6236 22491
rect 6184 22448 6236 22457
rect 7656 22448 7708 22500
rect 9588 22448 9640 22500
rect 9772 22448 9824 22500
rect 10968 22584 11020 22636
rect 10416 22559 10468 22568
rect 10416 22525 10425 22559
rect 10425 22525 10459 22559
rect 10459 22525 10468 22559
rect 10416 22516 10468 22525
rect 11060 22448 11112 22500
rect 11612 22559 11664 22568
rect 11612 22525 11621 22559
rect 11621 22525 11655 22559
rect 11655 22525 11664 22559
rect 11612 22516 11664 22525
rect 11520 22448 11572 22500
rect 11888 22559 11940 22568
rect 11888 22525 11897 22559
rect 11897 22525 11931 22559
rect 11931 22525 11940 22559
rect 11888 22516 11940 22525
rect 13176 22584 13228 22636
rect 12072 22516 12124 22568
rect 12256 22516 12308 22568
rect 12808 22491 12860 22500
rect 12808 22457 12817 22491
rect 12817 22457 12851 22491
rect 12851 22457 12860 22491
rect 12808 22448 12860 22457
rect 13268 22559 13320 22568
rect 13268 22525 13277 22559
rect 13277 22525 13311 22559
rect 13311 22525 13320 22559
rect 13268 22516 13320 22525
rect 13912 22652 13964 22704
rect 15752 22652 15804 22704
rect 13544 22627 13596 22636
rect 13544 22593 13553 22627
rect 13553 22593 13587 22627
rect 13587 22593 13596 22627
rect 13544 22584 13596 22593
rect 13820 22584 13872 22636
rect 16396 22720 16448 22772
rect 16764 22652 16816 22704
rect 16856 22652 16908 22704
rect 19064 22720 19116 22772
rect 18788 22652 18840 22704
rect 21456 22720 21508 22772
rect 13636 22516 13688 22568
rect 16028 22584 16080 22636
rect 13452 22448 13504 22500
rect 14648 22559 14700 22568
rect 14648 22525 14658 22559
rect 14658 22525 14692 22559
rect 14692 22525 14700 22559
rect 14648 22516 14700 22525
rect 14464 22491 14516 22500
rect 14464 22457 14473 22491
rect 14473 22457 14507 22491
rect 14507 22457 14516 22491
rect 14464 22448 14516 22457
rect 15108 22491 15160 22500
rect 15108 22457 15117 22491
rect 15117 22457 15151 22491
rect 15151 22457 15160 22491
rect 15108 22448 15160 22457
rect 16396 22516 16448 22568
rect 5080 22423 5132 22432
rect 5080 22389 5089 22423
rect 5089 22389 5123 22423
rect 5123 22389 5132 22423
rect 5080 22380 5132 22389
rect 5448 22380 5500 22432
rect 8484 22423 8536 22432
rect 8484 22389 8493 22423
rect 8493 22389 8527 22423
rect 8527 22389 8536 22423
rect 8484 22380 8536 22389
rect 9036 22423 9088 22432
rect 9036 22389 9045 22423
rect 9045 22389 9079 22423
rect 9079 22389 9088 22423
rect 9036 22380 9088 22389
rect 9864 22423 9916 22432
rect 9864 22389 9889 22423
rect 9889 22389 9916 22423
rect 9864 22380 9916 22389
rect 10048 22423 10100 22432
rect 10048 22389 10057 22423
rect 10057 22389 10091 22423
rect 10091 22389 10100 22423
rect 10048 22380 10100 22389
rect 11428 22380 11480 22432
rect 13360 22380 13412 22432
rect 16488 22491 16540 22500
rect 16488 22457 16497 22491
rect 16497 22457 16531 22491
rect 16531 22457 16540 22491
rect 16488 22448 16540 22457
rect 14924 22423 14976 22432
rect 14924 22389 14933 22423
rect 14933 22389 14967 22423
rect 14967 22389 14976 22423
rect 14924 22380 14976 22389
rect 15292 22423 15344 22432
rect 15292 22389 15317 22423
rect 15317 22389 15344 22423
rect 15292 22380 15344 22389
rect 15752 22380 15804 22432
rect 16304 22423 16356 22432
rect 16304 22389 16313 22423
rect 16313 22389 16347 22423
rect 16347 22389 16356 22423
rect 16304 22380 16356 22389
rect 16396 22380 16448 22432
rect 16856 22448 16908 22500
rect 17500 22491 17552 22500
rect 17500 22457 17509 22491
rect 17509 22457 17543 22491
rect 17543 22457 17552 22491
rect 17500 22448 17552 22457
rect 17592 22491 17644 22500
rect 17592 22457 17601 22491
rect 17601 22457 17635 22491
rect 17635 22457 17644 22491
rect 17592 22448 17644 22457
rect 17776 22491 17828 22500
rect 17776 22457 17785 22491
rect 17785 22457 17819 22491
rect 17819 22457 17828 22491
rect 17776 22448 17828 22457
rect 18696 22584 18748 22636
rect 19248 22627 19300 22636
rect 19248 22593 19257 22627
rect 19257 22593 19291 22627
rect 19291 22593 19300 22627
rect 19248 22584 19300 22593
rect 17960 22423 18012 22432
rect 17960 22389 17969 22423
rect 17969 22389 18003 22423
rect 18003 22389 18012 22423
rect 17960 22380 18012 22389
rect 19800 22559 19852 22568
rect 19800 22525 19809 22559
rect 19809 22525 19843 22559
rect 19843 22525 19852 22559
rect 19800 22516 19852 22525
rect 19984 22627 20036 22636
rect 19984 22593 19993 22627
rect 19993 22593 20027 22627
rect 20027 22593 20036 22627
rect 19984 22584 20036 22593
rect 20996 22584 21048 22636
rect 18420 22448 18472 22500
rect 18788 22448 18840 22500
rect 18880 22491 18932 22500
rect 18880 22457 18889 22491
rect 18889 22457 18923 22491
rect 18923 22457 18932 22491
rect 18880 22448 18932 22457
rect 18972 22448 19024 22500
rect 20536 22491 20588 22500
rect 20536 22457 20545 22491
rect 20545 22457 20579 22491
rect 20579 22457 20588 22491
rect 20536 22448 20588 22457
rect 21916 22720 21968 22772
rect 22008 22652 22060 22704
rect 22192 22448 22244 22500
rect 19064 22423 19116 22432
rect 19064 22389 19073 22423
rect 19073 22389 19107 22423
rect 19107 22389 19116 22423
rect 19064 22380 19116 22389
rect 21548 22380 21600 22432
rect 21640 22423 21692 22432
rect 21640 22389 21649 22423
rect 21649 22389 21683 22423
rect 21683 22389 21692 22423
rect 21640 22380 21692 22389
rect 4322 22278 4374 22330
rect 4386 22278 4438 22330
rect 4450 22278 4502 22330
rect 4514 22278 4566 22330
rect 4578 22278 4630 22330
rect 11612 22176 11664 22228
rect 7564 22108 7616 22160
rect 5632 22040 5684 22092
rect 6276 22083 6328 22092
rect 6276 22049 6285 22083
rect 6285 22049 6319 22083
rect 6319 22049 6328 22083
rect 6276 22040 6328 22049
rect 6920 22040 6972 22092
rect 8208 22040 8260 22092
rect 9220 22108 9272 22160
rect 10048 22108 10100 22160
rect 11244 22108 11296 22160
rect 9864 22040 9916 22092
rect 7380 21904 7432 21956
rect 7472 21947 7524 21956
rect 7472 21913 7481 21947
rect 7481 21913 7515 21947
rect 7515 21913 7524 21947
rect 7472 21904 7524 21913
rect 7656 21904 7708 21956
rect 8208 21904 8260 21956
rect 5264 21879 5316 21888
rect 5264 21845 5273 21879
rect 5273 21845 5307 21879
rect 5307 21845 5316 21879
rect 5264 21836 5316 21845
rect 6368 21836 6420 21888
rect 9220 21972 9272 22024
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 9680 21904 9732 21956
rect 10140 21904 10192 21956
rect 11152 22083 11204 22092
rect 11152 22049 11161 22083
rect 11161 22049 11195 22083
rect 11195 22049 11204 22083
rect 11152 22040 11204 22049
rect 11888 22108 11940 22160
rect 11796 22083 11848 22092
rect 11796 22049 11805 22083
rect 11805 22049 11839 22083
rect 11839 22049 11848 22083
rect 11796 22040 11848 22049
rect 12072 22083 12124 22092
rect 12072 22049 12081 22083
rect 12081 22049 12115 22083
rect 12115 22049 12124 22083
rect 12072 22040 12124 22049
rect 12808 22176 12860 22228
rect 14924 22176 14976 22228
rect 16304 22176 16356 22228
rect 10968 21972 11020 22024
rect 12716 22040 12768 22092
rect 13452 22040 13504 22092
rect 15568 22151 15620 22160
rect 15568 22117 15577 22151
rect 15577 22117 15611 22151
rect 15611 22117 15620 22151
rect 15568 22108 15620 22117
rect 17040 22108 17092 22160
rect 11336 21904 11388 21956
rect 13084 22015 13136 22024
rect 13084 21981 13093 22015
rect 13093 21981 13127 22015
rect 13127 21981 13136 22015
rect 13084 21972 13136 21981
rect 13820 22015 13872 22024
rect 13820 21981 13829 22015
rect 13829 21981 13863 22015
rect 13863 21981 13872 22015
rect 13820 21972 13872 21981
rect 14096 22083 14148 22092
rect 14096 22049 14105 22083
rect 14105 22049 14139 22083
rect 14139 22049 14148 22083
rect 14096 22040 14148 22049
rect 14648 22040 14700 22092
rect 15752 22083 15804 22092
rect 15752 22049 15761 22083
rect 15761 22049 15795 22083
rect 15795 22049 15804 22083
rect 15752 22040 15804 22049
rect 16120 22083 16172 22092
rect 16120 22049 16129 22083
rect 16129 22049 16163 22083
rect 16163 22049 16172 22083
rect 16120 22040 16172 22049
rect 16580 22083 16632 22092
rect 16580 22049 16589 22083
rect 16589 22049 16623 22083
rect 16623 22049 16632 22083
rect 16580 22040 16632 22049
rect 16764 22040 16816 22092
rect 17132 22040 17184 22092
rect 17408 22083 17460 22092
rect 17408 22049 17417 22083
rect 17417 22049 17451 22083
rect 17451 22049 17460 22083
rect 17408 22040 17460 22049
rect 18236 22176 18288 22228
rect 18788 22219 18840 22228
rect 18788 22185 18797 22219
rect 18797 22185 18831 22219
rect 18831 22185 18840 22219
rect 18788 22176 18840 22185
rect 21548 22176 21600 22228
rect 18420 22151 18472 22160
rect 18420 22117 18429 22151
rect 18429 22117 18463 22151
rect 18463 22117 18472 22151
rect 18420 22108 18472 22117
rect 21456 22108 21508 22160
rect 13636 21904 13688 21956
rect 15016 22015 15068 22024
rect 15016 21981 15025 22015
rect 15025 21981 15059 22015
rect 15059 21981 15068 22015
rect 15016 21972 15068 21981
rect 15476 21972 15528 22024
rect 16488 21972 16540 22024
rect 18972 22040 19024 22092
rect 19156 22040 19208 22092
rect 19708 22083 19760 22092
rect 19708 22049 19717 22083
rect 19717 22049 19751 22083
rect 19751 22049 19760 22083
rect 19708 22040 19760 22049
rect 19800 22040 19852 22092
rect 20996 22040 21048 22092
rect 17592 22015 17644 22024
rect 17592 21981 17601 22015
rect 17601 21981 17635 22015
rect 17635 21981 17644 22015
rect 17592 21972 17644 21981
rect 18144 21972 18196 22024
rect 19248 21972 19300 22024
rect 21548 22083 21600 22092
rect 21548 22049 21557 22083
rect 21557 22049 21591 22083
rect 21591 22049 21600 22083
rect 21548 22040 21600 22049
rect 21640 22083 21692 22092
rect 21640 22049 21649 22083
rect 21649 22049 21683 22083
rect 21683 22049 21692 22083
rect 21640 22040 21692 22049
rect 22560 22151 22612 22160
rect 22560 22117 22569 22151
rect 22569 22117 22603 22151
rect 22603 22117 22612 22151
rect 22560 22108 22612 22117
rect 15200 21904 15252 21956
rect 9404 21836 9456 21888
rect 12624 21836 12676 21888
rect 12992 21836 13044 21888
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 15476 21836 15528 21888
rect 17960 21836 18012 21888
rect 21180 21904 21232 21956
rect 21548 21904 21600 21956
rect 21824 21972 21876 22024
rect 22192 21972 22244 22024
rect 21916 21904 21968 21956
rect 19800 21836 19852 21888
rect 20628 21836 20680 21888
rect 21732 21879 21784 21888
rect 21732 21845 21741 21879
rect 21741 21845 21775 21879
rect 21775 21845 21784 21879
rect 21732 21836 21784 21845
rect 22100 21879 22152 21888
rect 22100 21845 22109 21879
rect 22109 21845 22143 21879
rect 22143 21845 22152 21879
rect 22100 21836 22152 21845
rect 3662 21734 3714 21786
rect 3726 21734 3778 21786
rect 3790 21734 3842 21786
rect 3854 21734 3906 21786
rect 3918 21734 3970 21786
rect 9036 21632 9088 21684
rect 9404 21632 9456 21684
rect 4712 21564 4764 21616
rect 5264 21607 5316 21616
rect 5264 21573 5273 21607
rect 5273 21573 5307 21607
rect 5307 21573 5316 21607
rect 5264 21564 5316 21573
rect 7564 21564 7616 21616
rect 9864 21564 9916 21616
rect 6184 21496 6236 21548
rect 6368 21496 6420 21548
rect 7196 21539 7248 21548
rect 7196 21505 7205 21539
rect 7205 21505 7239 21539
rect 7239 21505 7248 21539
rect 7196 21496 7248 21505
rect 7472 21496 7524 21548
rect 8484 21496 8536 21548
rect 5080 21360 5132 21412
rect 5264 21360 5316 21412
rect 6368 21403 6420 21412
rect 6368 21369 6377 21403
rect 6377 21369 6411 21403
rect 6411 21369 6420 21403
rect 6368 21360 6420 21369
rect 7748 21471 7800 21480
rect 7748 21437 7757 21471
rect 7757 21437 7791 21471
rect 7791 21437 7800 21471
rect 7748 21428 7800 21437
rect 8576 21428 8628 21480
rect 9220 21539 9272 21548
rect 9220 21505 9229 21539
rect 9229 21505 9263 21539
rect 9263 21505 9272 21539
rect 9220 21496 9272 21505
rect 9588 21428 9640 21480
rect 9772 21471 9824 21480
rect 9772 21437 9781 21471
rect 9781 21437 9815 21471
rect 9815 21437 9824 21471
rect 9772 21428 9824 21437
rect 7656 21360 7708 21412
rect 8116 21360 8168 21412
rect 8208 21360 8260 21412
rect 12164 21632 12216 21684
rect 13084 21632 13136 21684
rect 13452 21632 13504 21684
rect 10876 21607 10928 21616
rect 10876 21573 10885 21607
rect 10885 21573 10919 21607
rect 10919 21573 10928 21607
rect 10876 21564 10928 21573
rect 12624 21564 12676 21616
rect 10232 21428 10284 21480
rect 11980 21496 12032 21548
rect 12072 21539 12124 21548
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 12256 21496 12308 21548
rect 10784 21428 10836 21480
rect 5172 21292 5224 21344
rect 8484 21292 8536 21344
rect 9772 21292 9824 21344
rect 10784 21292 10836 21344
rect 12808 21428 12860 21480
rect 13268 21564 13320 21616
rect 13728 21564 13780 21616
rect 17224 21632 17276 21684
rect 17776 21632 17828 21684
rect 13544 21496 13596 21548
rect 14648 21539 14700 21548
rect 14648 21505 14657 21539
rect 14657 21505 14691 21539
rect 14691 21505 14700 21539
rect 14648 21496 14700 21505
rect 17408 21564 17460 21616
rect 19800 21632 19852 21684
rect 21456 21675 21508 21684
rect 21456 21641 21465 21675
rect 21465 21641 21499 21675
rect 21499 21641 21508 21675
rect 21456 21632 21508 21641
rect 18880 21564 18932 21616
rect 22192 21632 22244 21684
rect 17040 21496 17092 21548
rect 13360 21471 13412 21480
rect 13360 21437 13369 21471
rect 13369 21437 13403 21471
rect 13403 21437 13412 21471
rect 13360 21428 13412 21437
rect 12348 21360 12400 21412
rect 12716 21360 12768 21412
rect 14004 21471 14056 21480
rect 14004 21437 14013 21471
rect 14013 21437 14047 21471
rect 14047 21437 14056 21471
rect 14004 21428 14056 21437
rect 14464 21428 14516 21480
rect 14740 21471 14792 21480
rect 14740 21437 14749 21471
rect 14749 21437 14783 21471
rect 14783 21437 14792 21471
rect 14740 21428 14792 21437
rect 15936 21471 15988 21480
rect 15936 21437 15945 21471
rect 15945 21437 15979 21471
rect 15979 21437 15988 21471
rect 15936 21428 15988 21437
rect 16396 21428 16448 21480
rect 16120 21360 16172 21412
rect 17132 21471 17184 21480
rect 17132 21437 17141 21471
rect 17141 21437 17175 21471
rect 17175 21437 17184 21471
rect 17132 21428 17184 21437
rect 17316 21428 17368 21480
rect 17960 21471 18012 21480
rect 17960 21437 17969 21471
rect 17969 21437 18003 21471
rect 18003 21437 18012 21471
rect 17960 21428 18012 21437
rect 18420 21496 18472 21548
rect 18236 21471 18288 21480
rect 18236 21437 18245 21471
rect 18245 21437 18279 21471
rect 18279 21437 18288 21471
rect 18236 21428 18288 21437
rect 19064 21496 19116 21548
rect 19248 21539 19300 21548
rect 19248 21505 19257 21539
rect 19257 21505 19291 21539
rect 19291 21505 19300 21539
rect 19248 21496 19300 21505
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 17408 21360 17460 21412
rect 20536 21471 20588 21480
rect 20536 21437 20575 21471
rect 20575 21437 20588 21471
rect 20536 21428 20588 21437
rect 20720 21471 20772 21480
rect 20720 21437 20729 21471
rect 20729 21437 20763 21471
rect 20763 21437 20772 21471
rect 20720 21428 20772 21437
rect 20996 21471 21048 21480
rect 20996 21437 21005 21471
rect 21005 21437 21039 21471
rect 21039 21437 21048 21471
rect 20996 21428 21048 21437
rect 21088 21471 21140 21480
rect 21088 21437 21097 21471
rect 21097 21437 21131 21471
rect 21131 21437 21140 21471
rect 21088 21428 21140 21437
rect 21364 21428 21416 21480
rect 21180 21360 21232 21412
rect 12164 21335 12216 21344
rect 12164 21301 12173 21335
rect 12173 21301 12207 21335
rect 12207 21301 12216 21335
rect 12164 21292 12216 21301
rect 14096 21292 14148 21344
rect 14188 21335 14240 21344
rect 14188 21301 14197 21335
rect 14197 21301 14231 21335
rect 14231 21301 14240 21335
rect 14188 21292 14240 21301
rect 15292 21292 15344 21344
rect 17500 21335 17552 21344
rect 17500 21301 17509 21335
rect 17509 21301 17543 21335
rect 17543 21301 17552 21335
rect 17500 21292 17552 21301
rect 18880 21292 18932 21344
rect 20444 21292 20496 21344
rect 21916 21360 21968 21412
rect 22008 21292 22060 21344
rect 4322 21190 4374 21242
rect 4386 21190 4438 21242
rect 4450 21190 4502 21242
rect 4514 21190 4566 21242
rect 4578 21190 4630 21242
rect 5632 21088 5684 21140
rect 6368 21088 6420 21140
rect 5172 21020 5224 21072
rect 8116 21088 8168 21140
rect 5264 20952 5316 21004
rect 5632 20952 5684 21004
rect 7932 21020 7984 21072
rect 6920 20952 6972 21004
rect 7104 20952 7156 21004
rect 8208 20995 8260 21004
rect 8208 20961 8217 20995
rect 8217 20961 8251 20995
rect 8251 20961 8260 20995
rect 8208 20952 8260 20961
rect 9772 21088 9824 21140
rect 9404 21020 9456 21072
rect 9496 20995 9548 21004
rect 9496 20961 9505 20995
rect 9505 20961 9539 20995
rect 9539 20961 9548 20995
rect 9496 20952 9548 20961
rect 9680 20995 9732 21004
rect 9680 20961 9689 20995
rect 9689 20961 9723 20995
rect 9723 20961 9732 20995
rect 9680 20952 9732 20961
rect 9956 20952 10008 21004
rect 10784 21088 10836 21140
rect 11704 21088 11756 21140
rect 12348 21088 12400 21140
rect 14096 21131 14148 21140
rect 14096 21097 14105 21131
rect 14105 21097 14139 21131
rect 14139 21097 14148 21131
rect 14096 21088 14148 21097
rect 16488 21131 16540 21140
rect 16488 21097 16497 21131
rect 16497 21097 16531 21131
rect 16531 21097 16540 21131
rect 16488 21088 16540 21097
rect 17316 21131 17368 21140
rect 17316 21097 17325 21131
rect 17325 21097 17359 21131
rect 17359 21097 17368 21131
rect 17316 21088 17368 21097
rect 10324 20995 10376 21004
rect 10324 20961 10333 20995
rect 10333 20961 10367 20995
rect 10367 20961 10376 20995
rect 10324 20952 10376 20961
rect 10784 20995 10836 21004
rect 10784 20961 10793 20995
rect 10793 20961 10827 20995
rect 10827 20961 10836 20995
rect 10784 20952 10836 20961
rect 11060 20995 11112 21004
rect 11060 20961 11069 20995
rect 11069 20961 11103 20995
rect 11103 20961 11112 20995
rect 11060 20952 11112 20961
rect 11428 20995 11480 21004
rect 11428 20961 11437 20995
rect 11437 20961 11471 20995
rect 11471 20961 11480 20995
rect 11428 20952 11480 20961
rect 13176 20952 13228 21004
rect 13912 20995 13964 21004
rect 13912 20961 13921 20995
rect 13921 20961 13955 20995
rect 13955 20961 13964 20995
rect 13912 20952 13964 20961
rect 4620 20927 4672 20936
rect 4620 20893 4629 20927
rect 4629 20893 4663 20927
rect 4663 20893 4672 20927
rect 4620 20884 4672 20893
rect 5080 20884 5132 20936
rect 5356 20859 5408 20868
rect 5356 20825 5365 20859
rect 5365 20825 5399 20859
rect 5399 20825 5408 20859
rect 5356 20816 5408 20825
rect 11612 20884 11664 20936
rect 14924 21020 14976 21072
rect 15936 21020 15988 21072
rect 20996 21020 21048 21072
rect 15016 20952 15068 21004
rect 15476 20995 15528 21004
rect 15476 20961 15485 20995
rect 15485 20961 15519 20995
rect 15519 20961 15528 20995
rect 15476 20952 15528 20961
rect 16304 20995 16356 21004
rect 16304 20961 16313 20995
rect 16313 20961 16347 20995
rect 16347 20961 16356 20995
rect 16304 20952 16356 20961
rect 15752 20884 15804 20936
rect 17224 20995 17276 21004
rect 17224 20961 17233 20995
rect 17233 20961 17267 20995
rect 17267 20961 17276 20995
rect 17224 20952 17276 20961
rect 17592 20952 17644 21004
rect 20444 20995 20496 21004
rect 20444 20961 20453 20995
rect 20453 20961 20487 20995
rect 20487 20961 20496 20995
rect 20444 20952 20496 20961
rect 20536 20995 20588 21004
rect 20536 20961 20545 20995
rect 20545 20961 20579 20995
rect 20579 20961 20588 20995
rect 20536 20952 20588 20961
rect 20720 20995 20772 21004
rect 20720 20961 20733 20995
rect 20733 20961 20772 20995
rect 20720 20952 20772 20961
rect 21088 20952 21140 21004
rect 21732 20995 21784 21004
rect 21732 20961 21741 20995
rect 21741 20961 21775 20995
rect 21775 20961 21784 20995
rect 21732 20952 21784 20961
rect 5080 20748 5132 20800
rect 5448 20791 5500 20800
rect 5448 20757 5457 20791
rect 5457 20757 5491 20791
rect 5491 20757 5500 20791
rect 10324 20816 10376 20868
rect 15936 20816 15988 20868
rect 21548 20927 21600 20936
rect 21548 20893 21557 20927
rect 21557 20893 21591 20927
rect 21591 20893 21600 20927
rect 21548 20884 21600 20893
rect 22100 20859 22152 20868
rect 22100 20825 22109 20859
rect 22109 20825 22143 20859
rect 22143 20825 22152 20859
rect 22100 20816 22152 20825
rect 5448 20748 5500 20757
rect 6644 20748 6696 20800
rect 9128 20748 9180 20800
rect 9496 20748 9548 20800
rect 11152 20748 11204 20800
rect 11336 20748 11388 20800
rect 13728 20791 13780 20800
rect 13728 20757 13737 20791
rect 13737 20757 13771 20791
rect 13771 20757 13780 20791
rect 13728 20748 13780 20757
rect 20260 20748 20312 20800
rect 21272 20791 21324 20800
rect 21272 20757 21281 20791
rect 21281 20757 21315 20791
rect 21315 20757 21324 20791
rect 21272 20748 21324 20757
rect 21916 20791 21968 20800
rect 21916 20757 21925 20791
rect 21925 20757 21959 20791
rect 21959 20757 21968 20791
rect 21916 20748 21968 20757
rect 3662 20646 3714 20698
rect 3726 20646 3778 20698
rect 3790 20646 3842 20698
rect 3854 20646 3906 20698
rect 3918 20646 3970 20698
rect 5080 20587 5132 20596
rect 5080 20553 5089 20587
rect 5089 20553 5123 20587
rect 5123 20553 5132 20587
rect 5080 20544 5132 20553
rect 5448 20544 5500 20596
rect 6092 20544 6144 20596
rect 8668 20544 8720 20596
rect 10140 20544 10192 20596
rect 10784 20544 10836 20596
rect 13176 20544 13228 20596
rect 5172 20451 5224 20460
rect 5172 20417 5181 20451
rect 5181 20417 5215 20451
rect 5215 20417 5224 20451
rect 5172 20408 5224 20417
rect 5632 20451 5684 20460
rect 5632 20417 5641 20451
rect 5641 20417 5675 20451
rect 5675 20417 5684 20451
rect 5632 20408 5684 20417
rect 5908 20451 5960 20460
rect 5908 20417 5917 20451
rect 5917 20417 5951 20451
rect 5951 20417 5960 20451
rect 5908 20408 5960 20417
rect 5448 20340 5500 20392
rect 6000 20383 6052 20392
rect 6000 20349 6009 20383
rect 6009 20349 6043 20383
rect 6043 20349 6052 20383
rect 6000 20340 6052 20349
rect 6644 20383 6696 20392
rect 6644 20349 6653 20383
rect 6653 20349 6687 20383
rect 6687 20349 6696 20383
rect 6644 20340 6696 20349
rect 10876 20408 10928 20460
rect 12348 20408 12400 20460
rect 7104 20383 7156 20392
rect 7104 20349 7113 20383
rect 7113 20349 7147 20383
rect 7147 20349 7156 20383
rect 7104 20340 7156 20349
rect 7932 20340 7984 20392
rect 8576 20340 8628 20392
rect 8668 20383 8720 20392
rect 8668 20349 8677 20383
rect 8677 20349 8711 20383
rect 8711 20349 8720 20383
rect 8668 20340 8720 20349
rect 9680 20340 9732 20392
rect 10048 20340 10100 20392
rect 10968 20340 11020 20392
rect 12440 20340 12492 20392
rect 14648 20587 14700 20596
rect 14648 20553 14657 20587
rect 14657 20553 14691 20587
rect 14691 20553 14700 20587
rect 14648 20544 14700 20553
rect 15568 20476 15620 20528
rect 16304 20476 16356 20528
rect 14096 20408 14148 20460
rect 14372 20408 14424 20460
rect 16396 20408 16448 20460
rect 13728 20383 13780 20392
rect 13728 20349 13737 20383
rect 13737 20349 13771 20383
rect 13771 20349 13780 20383
rect 13728 20340 13780 20349
rect 14464 20383 14516 20392
rect 14464 20349 14473 20383
rect 14473 20349 14507 20383
rect 14507 20349 14516 20383
rect 14464 20340 14516 20349
rect 7380 20272 7432 20324
rect 17500 20340 17552 20392
rect 21548 20544 21600 20596
rect 22652 20476 22704 20528
rect 18328 20340 18380 20392
rect 18880 20383 18932 20392
rect 18880 20349 18889 20383
rect 18889 20349 18923 20383
rect 18923 20349 18932 20383
rect 18880 20340 18932 20349
rect 20536 20340 20588 20392
rect 5724 20204 5776 20256
rect 6368 20247 6420 20256
rect 6368 20213 6377 20247
rect 6377 20213 6411 20247
rect 6411 20213 6420 20247
rect 6368 20204 6420 20213
rect 6920 20204 6972 20256
rect 8944 20204 8996 20256
rect 13636 20204 13688 20256
rect 13820 20204 13872 20256
rect 17132 20204 17184 20256
rect 18144 20204 18196 20256
rect 18512 20204 18564 20256
rect 20444 20247 20496 20256
rect 20444 20213 20453 20247
rect 20453 20213 20487 20247
rect 20487 20213 20496 20247
rect 20444 20204 20496 20213
rect 20720 20383 20772 20392
rect 20720 20349 20729 20383
rect 20729 20349 20763 20383
rect 20763 20349 20772 20383
rect 20720 20340 20772 20349
rect 21088 20315 21140 20324
rect 21088 20281 21097 20315
rect 21097 20281 21131 20315
rect 21131 20281 21140 20315
rect 21088 20272 21140 20281
rect 21916 20340 21968 20392
rect 22192 20383 22244 20392
rect 22192 20349 22201 20383
rect 22201 20349 22235 20383
rect 22235 20349 22244 20383
rect 22192 20340 22244 20349
rect 21456 20247 21508 20256
rect 21456 20213 21465 20247
rect 21465 20213 21499 20247
rect 21499 20213 21508 20247
rect 21456 20204 21508 20213
rect 21640 20272 21692 20324
rect 22376 20247 22428 20256
rect 22376 20213 22385 20247
rect 22385 20213 22419 20247
rect 22419 20213 22428 20247
rect 22376 20204 22428 20213
rect 4322 20102 4374 20154
rect 4386 20102 4438 20154
rect 4450 20102 4502 20154
rect 4514 20102 4566 20154
rect 4578 20102 4630 20154
rect 7380 20043 7432 20052
rect 7380 20009 7389 20043
rect 7389 20009 7423 20043
rect 7423 20009 7432 20043
rect 7380 20000 7432 20009
rect 6000 19975 6052 19984
rect 6000 19941 6009 19975
rect 6009 19941 6043 19975
rect 6043 19941 6052 19975
rect 7932 20000 7984 20052
rect 6000 19932 6052 19941
rect 5540 19864 5592 19916
rect 6092 19864 6144 19916
rect 6920 19864 6972 19916
rect 7564 19907 7616 19916
rect 7564 19873 7573 19907
rect 7573 19873 7607 19907
rect 7607 19873 7616 19907
rect 7564 19864 7616 19873
rect 8576 19932 8628 19984
rect 13636 19975 13688 19984
rect 13636 19941 13645 19975
rect 13645 19941 13679 19975
rect 13679 19941 13688 19975
rect 13636 19932 13688 19941
rect 9772 19864 9824 19916
rect 10324 19907 10376 19916
rect 10324 19873 10333 19907
rect 10333 19873 10367 19907
rect 10367 19873 10376 19907
rect 10324 19864 10376 19873
rect 11060 19864 11112 19916
rect 12440 19907 12492 19916
rect 12440 19873 12449 19907
rect 12449 19873 12483 19907
rect 12483 19873 12492 19907
rect 12440 19864 12492 19873
rect 13176 19907 13228 19916
rect 13176 19873 13185 19907
rect 13185 19873 13219 19907
rect 13219 19873 13228 19907
rect 13176 19864 13228 19873
rect 13820 19907 13872 19916
rect 13820 19873 13829 19907
rect 13829 19873 13863 19907
rect 13863 19873 13872 19907
rect 13820 19864 13872 19873
rect 13912 19907 13964 19916
rect 13912 19873 13921 19907
rect 13921 19873 13955 19907
rect 13955 19873 13964 19907
rect 13912 19864 13964 19873
rect 14096 19864 14148 19916
rect 18144 20043 18196 20052
rect 18144 20009 18153 20043
rect 18153 20009 18187 20043
rect 18187 20009 18196 20043
rect 18144 20000 18196 20009
rect 18420 20000 18472 20052
rect 18788 20000 18840 20052
rect 19248 20043 19300 20052
rect 19248 20009 19275 20043
rect 19275 20009 19300 20043
rect 19248 20000 19300 20009
rect 20352 20000 20404 20052
rect 20720 20000 20772 20052
rect 21272 20043 21324 20052
rect 21272 20009 21281 20043
rect 21281 20009 21315 20043
rect 21315 20009 21324 20043
rect 21272 20000 21324 20009
rect 21456 20000 21508 20052
rect 16396 19864 16448 19916
rect 8300 19839 8352 19848
rect 8300 19805 8309 19839
rect 8309 19805 8343 19839
rect 8343 19805 8352 19839
rect 8300 19796 8352 19805
rect 11244 19839 11296 19848
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 12348 19839 12400 19848
rect 12348 19805 12357 19839
rect 12357 19805 12391 19839
rect 12391 19805 12400 19839
rect 12348 19796 12400 19805
rect 13728 19796 13780 19848
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 14832 19796 14884 19848
rect 6828 19728 6880 19780
rect 7748 19771 7800 19780
rect 7748 19737 7757 19771
rect 7757 19737 7791 19771
rect 7791 19737 7800 19771
rect 7748 19728 7800 19737
rect 9496 19728 9548 19780
rect 14740 19728 14792 19780
rect 17132 19907 17184 19916
rect 17132 19873 17141 19907
rect 17141 19873 17175 19907
rect 17175 19873 17184 19907
rect 17132 19864 17184 19873
rect 18420 19864 18472 19916
rect 18512 19907 18564 19916
rect 18512 19873 18521 19907
rect 18521 19873 18555 19907
rect 18555 19873 18564 19907
rect 18512 19864 18564 19873
rect 17960 19728 18012 19780
rect 10968 19660 11020 19712
rect 14372 19660 14424 19712
rect 15108 19660 15160 19712
rect 18788 19839 18840 19848
rect 18788 19805 18797 19839
rect 18797 19805 18831 19839
rect 18831 19805 18840 19839
rect 18788 19796 18840 19805
rect 19800 19907 19852 19916
rect 19800 19873 19809 19907
rect 19809 19873 19843 19907
rect 19843 19873 19852 19907
rect 19800 19864 19852 19873
rect 20260 19907 20312 19916
rect 20260 19873 20269 19907
rect 20269 19873 20303 19907
rect 20303 19873 20312 19907
rect 20260 19864 20312 19873
rect 20628 19907 20680 19916
rect 20628 19873 20637 19907
rect 20637 19873 20671 19907
rect 20671 19873 20680 19907
rect 20628 19864 20680 19873
rect 18328 19771 18380 19780
rect 18328 19737 18337 19771
rect 18337 19737 18371 19771
rect 18371 19737 18380 19771
rect 18328 19728 18380 19737
rect 19064 19703 19116 19712
rect 19064 19669 19073 19703
rect 19073 19669 19107 19703
rect 19107 19669 19116 19703
rect 19064 19660 19116 19669
rect 20628 19728 20680 19780
rect 21088 19907 21140 19916
rect 21088 19873 21097 19907
rect 21097 19873 21131 19907
rect 21131 19873 21140 19907
rect 21088 19864 21140 19873
rect 22284 19907 22336 19916
rect 22284 19873 22293 19907
rect 22293 19873 22327 19907
rect 22327 19873 22336 19907
rect 22284 19864 22336 19873
rect 22376 19907 22428 19916
rect 22376 19873 22385 19907
rect 22385 19873 22419 19907
rect 22419 19873 22428 19907
rect 22376 19864 22428 19873
rect 20996 19796 21048 19848
rect 21732 19839 21784 19848
rect 21732 19805 21741 19839
rect 21741 19805 21775 19839
rect 21775 19805 21784 19839
rect 21732 19796 21784 19805
rect 20260 19703 20312 19712
rect 20260 19669 20269 19703
rect 20269 19669 20303 19703
rect 20303 19669 20312 19703
rect 20260 19660 20312 19669
rect 22468 19660 22520 19712
rect 22652 19703 22704 19712
rect 22652 19669 22661 19703
rect 22661 19669 22695 19703
rect 22695 19669 22704 19703
rect 22652 19660 22704 19669
rect 22744 19660 22796 19712
rect 3662 19558 3714 19610
rect 3726 19558 3778 19610
rect 3790 19558 3842 19610
rect 3854 19558 3906 19610
rect 3918 19558 3970 19610
rect 5632 19499 5684 19508
rect 5632 19465 5641 19499
rect 5641 19465 5675 19499
rect 5675 19465 5684 19499
rect 5632 19456 5684 19465
rect 7564 19456 7616 19508
rect 7748 19363 7800 19372
rect 7748 19329 7757 19363
rect 7757 19329 7791 19363
rect 7791 19329 7800 19363
rect 7748 19320 7800 19329
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 6920 19252 6972 19304
rect 4712 19184 4764 19236
rect 5448 19227 5500 19236
rect 5448 19193 5457 19227
rect 5457 19193 5491 19227
rect 5491 19193 5500 19227
rect 5448 19184 5500 19193
rect 7564 19184 7616 19236
rect 8668 19295 8720 19304
rect 8668 19261 8677 19295
rect 8677 19261 8711 19295
rect 8711 19261 8720 19295
rect 8668 19252 8720 19261
rect 9404 19252 9456 19304
rect 13636 19388 13688 19440
rect 10968 19252 11020 19304
rect 11980 19295 12032 19304
rect 11980 19261 11989 19295
rect 11989 19261 12023 19295
rect 12023 19261 12032 19295
rect 11980 19252 12032 19261
rect 5264 19116 5316 19168
rect 7288 19116 7340 19168
rect 9588 19116 9640 19168
rect 11060 19184 11112 19236
rect 12348 19184 12400 19236
rect 13728 19252 13780 19304
rect 13820 19295 13872 19304
rect 13820 19261 13829 19295
rect 13829 19261 13863 19295
rect 13863 19261 13872 19295
rect 13820 19252 13872 19261
rect 14096 19295 14148 19304
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 14280 19295 14332 19304
rect 14280 19261 14293 19295
rect 14293 19261 14332 19295
rect 14280 19252 14332 19261
rect 14556 19295 14608 19304
rect 14556 19261 14565 19295
rect 14565 19261 14599 19295
rect 14599 19261 14608 19295
rect 14556 19252 14608 19261
rect 14740 19295 14792 19304
rect 14740 19261 14749 19295
rect 14749 19261 14783 19295
rect 14783 19261 14792 19295
rect 14740 19252 14792 19261
rect 18696 19456 18748 19508
rect 18880 19456 18932 19508
rect 22560 19456 22612 19508
rect 15476 19363 15528 19372
rect 15476 19329 15485 19363
rect 15485 19329 15519 19363
rect 15519 19329 15528 19363
rect 15476 19320 15528 19329
rect 15476 19184 15528 19236
rect 16304 19295 16356 19304
rect 16304 19261 16313 19295
rect 16313 19261 16347 19295
rect 16347 19261 16356 19295
rect 16304 19252 16356 19261
rect 16396 19295 16448 19304
rect 16396 19261 16405 19295
rect 16405 19261 16439 19295
rect 16439 19261 16448 19295
rect 16396 19252 16448 19261
rect 18328 19388 18380 19440
rect 17960 19295 18012 19304
rect 17960 19261 17969 19295
rect 17969 19261 18003 19295
rect 18003 19261 18012 19295
rect 17960 19252 18012 19261
rect 20260 19388 20312 19440
rect 20444 19388 20496 19440
rect 19064 19252 19116 19304
rect 20260 19295 20312 19304
rect 20260 19261 20269 19295
rect 20269 19261 20303 19295
rect 20303 19261 20312 19295
rect 20260 19252 20312 19261
rect 19340 19184 19392 19236
rect 20444 19295 20496 19304
rect 20444 19261 20453 19295
rect 20453 19261 20487 19295
rect 20487 19261 20496 19295
rect 20444 19252 20496 19261
rect 20628 19295 20680 19304
rect 10140 19116 10192 19168
rect 14464 19159 14516 19168
rect 14464 19125 14473 19159
rect 14473 19125 14507 19159
rect 14507 19125 14516 19159
rect 14464 19116 14516 19125
rect 14740 19116 14792 19168
rect 15384 19116 15436 19168
rect 18236 19159 18288 19168
rect 18236 19125 18245 19159
rect 18245 19125 18279 19159
rect 18279 19125 18288 19159
rect 18236 19116 18288 19125
rect 18512 19116 18564 19168
rect 19984 19159 20036 19168
rect 19984 19125 19993 19159
rect 19993 19125 20027 19159
rect 20027 19125 20036 19159
rect 19984 19116 20036 19125
rect 20168 19116 20220 19168
rect 20628 19261 20637 19295
rect 20637 19261 20671 19295
rect 20671 19261 20680 19295
rect 20628 19252 20680 19261
rect 21088 19295 21140 19304
rect 21088 19261 21100 19295
rect 21100 19261 21134 19295
rect 21134 19261 21140 19295
rect 21088 19252 21140 19261
rect 22468 19295 22520 19304
rect 22468 19261 22486 19295
rect 22486 19261 22520 19295
rect 22468 19252 22520 19261
rect 22836 19252 22888 19304
rect 21732 19184 21784 19236
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 22284 19116 22336 19168
rect 4322 19014 4374 19066
rect 4386 19014 4438 19066
rect 4450 19014 4502 19066
rect 4514 19014 4566 19066
rect 4578 19014 4630 19066
rect 6000 18912 6052 18964
rect 7564 18912 7616 18964
rect 8300 18955 8352 18964
rect 8300 18921 8309 18955
rect 8309 18921 8343 18955
rect 8343 18921 8352 18955
rect 8300 18912 8352 18921
rect 5448 18776 5500 18828
rect 5540 18708 5592 18760
rect 5264 18640 5316 18692
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 6828 18819 6880 18828
rect 6828 18785 6837 18819
rect 6837 18785 6871 18819
rect 6871 18785 6880 18819
rect 6828 18776 6880 18785
rect 7196 18776 7248 18828
rect 8392 18844 8444 18896
rect 11244 18912 11296 18964
rect 14464 18912 14516 18964
rect 10048 18887 10100 18896
rect 10048 18853 10057 18887
rect 10057 18853 10091 18887
rect 10091 18853 10100 18887
rect 10048 18844 10100 18853
rect 12072 18887 12124 18896
rect 12072 18853 12081 18887
rect 12081 18853 12115 18887
rect 12115 18853 12124 18887
rect 12072 18844 12124 18853
rect 7472 18819 7524 18828
rect 7472 18785 7481 18819
rect 7481 18785 7515 18819
rect 7515 18785 7524 18819
rect 7472 18776 7524 18785
rect 8852 18819 8904 18828
rect 8852 18785 8861 18819
rect 8861 18785 8895 18819
rect 8895 18785 8904 18819
rect 8852 18776 8904 18785
rect 8944 18819 8996 18828
rect 8944 18785 8953 18819
rect 8953 18785 8987 18819
rect 8987 18785 8996 18819
rect 8944 18776 8996 18785
rect 9404 18776 9456 18828
rect 7748 18708 7800 18760
rect 8760 18708 8812 18760
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 10600 18819 10652 18828
rect 10600 18785 10609 18819
rect 10609 18785 10643 18819
rect 10643 18785 10652 18819
rect 10600 18776 10652 18785
rect 10968 18819 11020 18828
rect 10968 18785 10977 18819
rect 10977 18785 11011 18819
rect 11011 18785 11020 18819
rect 10968 18776 11020 18785
rect 11336 18819 11388 18828
rect 11336 18785 11345 18819
rect 11345 18785 11379 18819
rect 11379 18785 11388 18819
rect 11336 18776 11388 18785
rect 11704 18776 11756 18828
rect 13636 18819 13688 18828
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 13728 18819 13780 18828
rect 13728 18785 13737 18819
rect 13737 18785 13771 18819
rect 13771 18785 13780 18819
rect 13728 18776 13780 18785
rect 14372 18776 14424 18828
rect 14648 18844 14700 18896
rect 14740 18819 14792 18828
rect 14740 18785 14749 18819
rect 14749 18785 14783 18819
rect 14783 18785 14792 18819
rect 14740 18776 14792 18785
rect 15108 18776 15160 18828
rect 15384 18776 15436 18828
rect 20536 18912 20588 18964
rect 22376 18912 22428 18964
rect 22560 18912 22612 18964
rect 16396 18844 16448 18896
rect 18236 18844 18288 18896
rect 18696 18819 18748 18828
rect 18696 18785 18705 18819
rect 18705 18785 18739 18819
rect 18739 18785 18748 18819
rect 18696 18776 18748 18785
rect 19984 18844 20036 18896
rect 21272 18844 21324 18896
rect 9496 18708 9548 18717
rect 10324 18708 10376 18760
rect 11980 18708 12032 18760
rect 13820 18640 13872 18692
rect 6736 18572 6788 18624
rect 9404 18572 9456 18624
rect 10048 18572 10100 18624
rect 11612 18572 11664 18624
rect 16304 18708 16356 18760
rect 18512 18708 18564 18760
rect 18880 18708 18932 18760
rect 21916 18776 21968 18828
rect 22928 18819 22980 18828
rect 22928 18785 22937 18819
rect 22937 18785 22971 18819
rect 22971 18785 22980 18819
rect 22928 18776 22980 18785
rect 19524 18751 19576 18760
rect 19524 18717 19533 18751
rect 19533 18717 19567 18751
rect 19567 18717 19576 18751
rect 19524 18708 19576 18717
rect 14464 18683 14516 18692
rect 14464 18649 14473 18683
rect 14473 18649 14507 18683
rect 14507 18649 14516 18683
rect 14464 18640 14516 18649
rect 16120 18683 16172 18692
rect 16120 18649 16129 18683
rect 16129 18649 16163 18683
rect 16163 18649 16172 18683
rect 16120 18640 16172 18649
rect 15016 18615 15068 18624
rect 15016 18581 15025 18615
rect 15025 18581 15059 18615
rect 15059 18581 15068 18615
rect 15016 18572 15068 18581
rect 15108 18572 15160 18624
rect 18512 18615 18564 18624
rect 18512 18581 18521 18615
rect 18521 18581 18555 18615
rect 18555 18581 18564 18615
rect 18512 18572 18564 18581
rect 18696 18572 18748 18624
rect 18788 18615 18840 18624
rect 18788 18581 18797 18615
rect 18797 18581 18831 18615
rect 18831 18581 18840 18615
rect 18788 18572 18840 18581
rect 20904 18615 20956 18624
rect 20904 18581 20913 18615
rect 20913 18581 20947 18615
rect 20947 18581 20956 18615
rect 20904 18572 20956 18581
rect 21548 18572 21600 18624
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 5632 18368 5684 18420
rect 6828 18368 6880 18420
rect 8760 18411 8812 18420
rect 8760 18377 8769 18411
rect 8769 18377 8803 18411
rect 8803 18377 8812 18411
rect 8760 18368 8812 18377
rect 10416 18368 10468 18420
rect 11336 18368 11388 18420
rect 5264 18275 5316 18284
rect 5264 18241 5273 18275
rect 5273 18241 5307 18275
rect 5307 18241 5316 18275
rect 5264 18232 5316 18241
rect 6736 18275 6788 18284
rect 6736 18241 6745 18275
rect 6745 18241 6779 18275
rect 6779 18241 6788 18275
rect 6736 18232 6788 18241
rect 4804 18164 4856 18216
rect 5448 18164 5500 18216
rect 6000 18164 6052 18216
rect 7012 18232 7064 18284
rect 7196 18275 7248 18284
rect 7196 18241 7205 18275
rect 7205 18241 7239 18275
rect 7239 18241 7248 18275
rect 7196 18232 7248 18241
rect 7288 18275 7340 18284
rect 7288 18241 7297 18275
rect 7297 18241 7331 18275
rect 7331 18241 7340 18275
rect 7288 18232 7340 18241
rect 4712 18096 4764 18148
rect 5356 18096 5408 18148
rect 6368 18096 6420 18148
rect 7748 18164 7800 18216
rect 8024 18232 8076 18284
rect 10600 18300 10652 18352
rect 10968 18300 11020 18352
rect 11704 18300 11756 18352
rect 14556 18368 14608 18420
rect 19800 18368 19852 18420
rect 20444 18368 20496 18420
rect 21640 18368 21692 18420
rect 13268 18300 13320 18352
rect 14372 18300 14424 18352
rect 8116 18207 8168 18216
rect 8116 18173 8125 18207
rect 8125 18173 8159 18207
rect 8159 18173 8168 18207
rect 8116 18164 8168 18173
rect 8392 18207 8444 18216
rect 8392 18173 8401 18207
rect 8401 18173 8435 18207
rect 8435 18173 8444 18207
rect 8392 18164 8444 18173
rect 8852 18164 8904 18216
rect 9036 18164 9088 18216
rect 9772 18207 9824 18216
rect 9772 18173 9781 18207
rect 9781 18173 9815 18207
rect 9815 18173 9824 18207
rect 9772 18164 9824 18173
rect 10324 18164 10376 18216
rect 11612 18207 11664 18216
rect 11612 18173 11621 18207
rect 11621 18173 11655 18207
rect 11655 18173 11664 18207
rect 11612 18164 11664 18173
rect 15016 18232 15068 18284
rect 11980 18207 12032 18216
rect 11980 18173 11989 18207
rect 11989 18173 12023 18207
rect 12023 18173 12032 18207
rect 11980 18164 12032 18173
rect 11060 18096 11112 18148
rect 11888 18139 11940 18148
rect 11888 18105 11897 18139
rect 11897 18105 11931 18139
rect 11931 18105 11940 18139
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 14924 18164 14976 18216
rect 18604 18300 18656 18352
rect 15752 18232 15804 18284
rect 15384 18207 15436 18216
rect 15384 18173 15393 18207
rect 15393 18173 15427 18207
rect 15427 18173 15436 18207
rect 15384 18164 15436 18173
rect 15660 18164 15712 18216
rect 16120 18164 16172 18216
rect 17500 18207 17552 18216
rect 17500 18173 17509 18207
rect 17509 18173 17543 18207
rect 17543 18173 17552 18207
rect 17500 18164 17552 18173
rect 17684 18207 17736 18216
rect 17684 18173 17693 18207
rect 17693 18173 17727 18207
rect 17727 18173 17736 18207
rect 17684 18164 17736 18173
rect 18696 18232 18748 18284
rect 18972 18275 19024 18284
rect 18972 18241 18981 18275
rect 18981 18241 19015 18275
rect 19015 18241 19024 18275
rect 18972 18232 19024 18241
rect 20904 18232 20956 18284
rect 11888 18096 11940 18105
rect 15476 18096 15528 18148
rect 17592 18096 17644 18148
rect 18604 18164 18656 18216
rect 18788 18164 18840 18216
rect 18880 18207 18932 18216
rect 18880 18173 18889 18207
rect 18889 18173 18923 18207
rect 18923 18173 18932 18207
rect 18880 18164 18932 18173
rect 19340 18164 19392 18216
rect 20536 18207 20588 18216
rect 20536 18173 20545 18207
rect 20545 18173 20579 18207
rect 20579 18173 20588 18207
rect 20536 18164 20588 18173
rect 21272 18207 21324 18216
rect 21272 18173 21281 18207
rect 21281 18173 21315 18207
rect 21315 18173 21324 18207
rect 21272 18164 21324 18173
rect 21640 18207 21692 18216
rect 21640 18173 21649 18207
rect 21649 18173 21683 18207
rect 21683 18173 21692 18207
rect 21640 18164 21692 18173
rect 21548 18139 21600 18148
rect 21548 18105 21557 18139
rect 21557 18105 21591 18139
rect 21591 18105 21600 18139
rect 21548 18096 21600 18105
rect 6276 18028 6328 18080
rect 6552 18071 6604 18080
rect 6552 18037 6561 18071
rect 6561 18037 6595 18071
rect 6595 18037 6604 18071
rect 6552 18028 6604 18037
rect 7104 18028 7156 18080
rect 8116 18028 8168 18080
rect 9864 18028 9916 18080
rect 15568 18071 15620 18080
rect 15568 18037 15577 18071
rect 15577 18037 15611 18071
rect 15611 18037 15620 18071
rect 15568 18028 15620 18037
rect 16764 18028 16816 18080
rect 16856 18071 16908 18080
rect 16856 18037 16865 18071
rect 16865 18037 16899 18071
rect 16899 18037 16908 18071
rect 16856 18028 16908 18037
rect 18696 18071 18748 18080
rect 18696 18037 18705 18071
rect 18705 18037 18739 18071
rect 18739 18037 18748 18071
rect 18696 18028 18748 18037
rect 21916 18028 21968 18080
rect 22376 18028 22428 18080
rect 22928 18028 22980 18080
rect 4322 17926 4374 17978
rect 4386 17926 4438 17978
rect 4450 17926 4502 17978
rect 4514 17926 4566 17978
rect 4578 17926 4630 17978
rect 5172 17824 5224 17876
rect 5540 17824 5592 17876
rect 4804 17799 4856 17808
rect 4804 17765 4813 17799
rect 4813 17765 4847 17799
rect 4847 17765 4856 17799
rect 4804 17756 4856 17765
rect 5264 17799 5316 17808
rect 5264 17765 5273 17799
rect 5273 17765 5307 17799
rect 5307 17765 5316 17799
rect 5264 17756 5316 17765
rect 10324 17867 10376 17876
rect 10324 17833 10333 17867
rect 10333 17833 10367 17867
rect 10367 17833 10376 17867
rect 10324 17824 10376 17833
rect 5356 17731 5408 17740
rect 5356 17697 5365 17731
rect 5365 17697 5399 17731
rect 5399 17697 5408 17731
rect 5356 17688 5408 17697
rect 5632 17688 5684 17740
rect 5540 17620 5592 17672
rect 6276 17688 6328 17740
rect 6552 17688 6604 17740
rect 10784 17756 10836 17808
rect 14464 17824 14516 17876
rect 16028 17824 16080 17876
rect 17684 17824 17736 17876
rect 6000 17663 6052 17672
rect 6000 17629 6009 17663
rect 6009 17629 6043 17663
rect 6043 17629 6052 17663
rect 6000 17620 6052 17629
rect 7012 17620 7064 17672
rect 7196 17620 7248 17672
rect 9680 17688 9732 17740
rect 10232 17688 10284 17740
rect 10968 17731 11020 17740
rect 10968 17697 10977 17731
rect 10977 17697 11011 17731
rect 11011 17697 11020 17731
rect 10968 17688 11020 17697
rect 12072 17688 12124 17740
rect 12532 17688 12584 17740
rect 16120 17799 16172 17808
rect 8576 17620 8628 17672
rect 10140 17620 10192 17672
rect 12348 17663 12400 17672
rect 12348 17629 12357 17663
rect 12357 17629 12391 17663
rect 12391 17629 12400 17663
rect 12348 17620 12400 17629
rect 13268 17663 13320 17672
rect 13268 17629 13277 17663
rect 13277 17629 13311 17663
rect 13311 17629 13320 17663
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 15752 17731 15804 17740
rect 15752 17697 15761 17731
rect 15761 17697 15795 17731
rect 15795 17697 15804 17731
rect 15752 17688 15804 17697
rect 13268 17620 13320 17629
rect 16120 17765 16129 17799
rect 16129 17765 16163 17799
rect 16163 17765 16172 17799
rect 16120 17756 16172 17765
rect 17132 17756 17184 17808
rect 16856 17688 16908 17740
rect 17408 17688 17460 17740
rect 16304 17620 16356 17672
rect 16488 17620 16540 17672
rect 17316 17620 17368 17672
rect 18236 17688 18288 17740
rect 18512 17799 18564 17808
rect 18512 17765 18521 17799
rect 18521 17765 18555 17799
rect 18555 17765 18564 17799
rect 18512 17756 18564 17765
rect 21548 17824 21600 17876
rect 23020 17799 23072 17808
rect 23020 17765 23029 17799
rect 23029 17765 23063 17799
rect 23063 17765 23072 17799
rect 23020 17756 23072 17765
rect 18144 17620 18196 17672
rect 5448 17484 5500 17536
rect 6460 17484 6512 17536
rect 8852 17484 8904 17536
rect 10048 17484 10100 17536
rect 16028 17552 16080 17604
rect 16212 17484 16264 17536
rect 17592 17552 17644 17604
rect 18328 17552 18380 17604
rect 18052 17484 18104 17536
rect 18696 17731 18748 17740
rect 18696 17697 18705 17731
rect 18705 17697 18739 17731
rect 18739 17697 18748 17731
rect 18696 17688 18748 17697
rect 19524 17688 19576 17740
rect 21272 17688 21324 17740
rect 21824 17731 21876 17740
rect 21824 17697 21833 17731
rect 21833 17697 21867 17731
rect 21867 17697 21876 17731
rect 21824 17688 21876 17697
rect 21916 17731 21968 17740
rect 21916 17697 21925 17731
rect 21925 17697 21959 17731
rect 21959 17697 21968 17731
rect 21916 17688 21968 17697
rect 22376 17731 22428 17740
rect 22376 17697 22385 17731
rect 22385 17697 22419 17731
rect 22419 17697 22428 17731
rect 22376 17688 22428 17697
rect 22560 17731 22612 17740
rect 22560 17697 22569 17731
rect 22569 17697 22603 17731
rect 22603 17697 22612 17731
rect 22560 17688 22612 17697
rect 20812 17620 20864 17672
rect 22192 17620 22244 17672
rect 18696 17552 18748 17604
rect 22100 17552 22152 17604
rect 22836 17620 22888 17672
rect 19432 17484 19484 17536
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 5264 17119 5316 17128
rect 5264 17085 5273 17119
rect 5273 17085 5307 17119
rect 5307 17085 5316 17119
rect 5264 17076 5316 17085
rect 5356 17119 5408 17128
rect 5356 17085 5365 17119
rect 5365 17085 5399 17119
rect 5399 17085 5408 17119
rect 5356 17076 5408 17085
rect 5448 17119 5500 17128
rect 5448 17085 5457 17119
rect 5457 17085 5491 17119
rect 5491 17085 5500 17119
rect 5448 17076 5500 17085
rect 6000 17280 6052 17332
rect 6920 17280 6972 17332
rect 9496 17280 9548 17332
rect 5908 17212 5960 17264
rect 6368 17212 6420 17264
rect 9036 17212 9088 17264
rect 9864 17212 9916 17264
rect 5816 17051 5868 17060
rect 5816 17017 5825 17051
rect 5825 17017 5859 17051
rect 5859 17017 5868 17051
rect 5816 17008 5868 17017
rect 5172 16940 5224 16992
rect 6368 17119 6420 17128
rect 6368 17085 6377 17119
rect 6377 17085 6411 17119
rect 6411 17085 6420 17119
rect 6368 17076 6420 17085
rect 6460 17119 6512 17128
rect 6460 17085 6469 17119
rect 6469 17085 6503 17119
rect 6503 17085 6512 17119
rect 6460 17076 6512 17085
rect 6552 17076 6604 17128
rect 7012 17119 7064 17128
rect 7012 17085 7021 17119
rect 7021 17085 7055 17119
rect 7055 17085 7064 17119
rect 7012 17076 7064 17085
rect 8852 17119 8904 17128
rect 8852 17085 8861 17119
rect 8861 17085 8895 17119
rect 8895 17085 8904 17119
rect 8852 17076 8904 17085
rect 9312 17076 9364 17128
rect 9680 17119 9732 17128
rect 9680 17085 9689 17119
rect 9689 17085 9723 17119
rect 9723 17085 9732 17119
rect 9680 17076 9732 17085
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 10968 17280 11020 17332
rect 12348 17280 12400 17332
rect 15016 17323 15068 17332
rect 15016 17289 15025 17323
rect 15025 17289 15059 17323
rect 15059 17289 15068 17323
rect 15016 17280 15068 17289
rect 15384 17212 15436 17264
rect 17132 17323 17184 17332
rect 17132 17289 17141 17323
rect 17141 17289 17175 17323
rect 17175 17289 17184 17323
rect 17132 17280 17184 17289
rect 17408 17323 17460 17332
rect 17408 17289 17417 17323
rect 17417 17289 17451 17323
rect 17451 17289 17460 17323
rect 17408 17280 17460 17289
rect 17684 17323 17736 17332
rect 17684 17289 17693 17323
rect 17693 17289 17727 17323
rect 17727 17289 17736 17323
rect 17684 17280 17736 17289
rect 18144 17323 18196 17332
rect 18144 17289 18153 17323
rect 18153 17289 18187 17323
rect 18187 17289 18196 17323
rect 18144 17280 18196 17289
rect 18972 17280 19024 17332
rect 16488 17212 16540 17264
rect 16948 17255 17000 17264
rect 16948 17221 16957 17255
rect 16957 17221 16991 17255
rect 16991 17221 17000 17255
rect 16948 17212 17000 17221
rect 15568 17187 15620 17196
rect 10416 17076 10468 17128
rect 10784 17119 10836 17128
rect 10784 17085 10793 17119
rect 10793 17085 10827 17119
rect 10827 17085 10836 17119
rect 10784 17076 10836 17085
rect 15568 17153 15577 17187
rect 15577 17153 15611 17187
rect 15611 17153 15620 17187
rect 15568 17144 15620 17153
rect 16304 17187 16356 17196
rect 16304 17153 16313 17187
rect 16313 17153 16347 17187
rect 16347 17153 16356 17187
rect 16304 17144 16356 17153
rect 16856 17144 16908 17196
rect 17500 17144 17552 17196
rect 14648 17119 14700 17128
rect 14648 17085 14657 17119
rect 14657 17085 14691 17119
rect 14691 17085 14700 17119
rect 14648 17076 14700 17085
rect 14464 17008 14516 17060
rect 16120 17076 16172 17128
rect 16672 17119 16724 17128
rect 16672 17085 16681 17119
rect 16681 17085 16715 17119
rect 16715 17085 16724 17119
rect 16672 17076 16724 17085
rect 16764 17076 16816 17128
rect 15200 17051 15252 17060
rect 15200 17017 15209 17051
rect 15209 17017 15243 17051
rect 15243 17017 15252 17051
rect 15200 17008 15252 17017
rect 16856 17008 16908 17060
rect 17132 17008 17184 17060
rect 6092 16983 6144 16992
rect 6092 16949 6101 16983
rect 6101 16949 6135 16983
rect 6135 16949 6144 16983
rect 6092 16940 6144 16949
rect 9772 16940 9824 16992
rect 9956 16983 10008 16992
rect 9956 16949 9965 16983
rect 9965 16949 9999 16983
rect 9999 16949 10008 16983
rect 9956 16940 10008 16949
rect 14648 16940 14700 16992
rect 16212 16940 16264 16992
rect 16764 16983 16816 16992
rect 16764 16949 16773 16983
rect 16773 16949 16807 16983
rect 16807 16949 16816 16983
rect 17592 17119 17644 17128
rect 17592 17085 17601 17119
rect 17601 17085 17635 17119
rect 17635 17085 17644 17119
rect 17592 17076 17644 17085
rect 18052 17144 18104 17196
rect 18420 17076 18472 17128
rect 18604 17076 18656 17128
rect 18696 17119 18748 17128
rect 18696 17085 18705 17119
rect 18705 17085 18739 17119
rect 18739 17085 18748 17119
rect 18696 17076 18748 17085
rect 19524 17076 19576 17128
rect 22100 17280 22152 17332
rect 22192 17280 22244 17332
rect 17408 17008 17460 17060
rect 19984 17008 20036 17060
rect 21640 17076 21692 17128
rect 22192 17076 22244 17128
rect 21272 17008 21324 17060
rect 16764 16940 16816 16949
rect 17500 16940 17552 16992
rect 19340 16940 19392 16992
rect 20076 16983 20128 16992
rect 20076 16949 20085 16983
rect 20085 16949 20119 16983
rect 20119 16949 20128 16983
rect 20076 16940 20128 16949
rect 21732 16940 21784 16992
rect 4322 16838 4374 16890
rect 4386 16838 4438 16890
rect 4450 16838 4502 16890
rect 4514 16838 4566 16890
rect 4578 16838 4630 16890
rect 4896 16736 4948 16788
rect 9496 16779 9548 16788
rect 9496 16745 9505 16779
rect 9505 16745 9539 16779
rect 9539 16745 9548 16779
rect 9496 16736 9548 16745
rect 9956 16736 10008 16788
rect 14464 16779 14516 16788
rect 14464 16745 14473 16779
rect 14473 16745 14507 16779
rect 14507 16745 14516 16779
rect 14464 16736 14516 16745
rect 16672 16736 16724 16788
rect 18236 16736 18288 16788
rect 19340 16736 19392 16788
rect 5448 16668 5500 16720
rect 4712 16643 4764 16652
rect 4712 16609 4721 16643
rect 4721 16609 4755 16643
rect 4755 16609 4764 16643
rect 4712 16600 4764 16609
rect 4804 16600 4856 16652
rect 5908 16600 5960 16652
rect 5540 16532 5592 16584
rect 5816 16532 5868 16584
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 7472 16668 7524 16720
rect 8576 16668 8628 16720
rect 7104 16643 7156 16652
rect 7104 16609 7113 16643
rect 7113 16609 7147 16643
rect 7147 16609 7156 16643
rect 7104 16600 7156 16609
rect 9312 16643 9364 16652
rect 9312 16609 9321 16643
rect 9321 16609 9355 16643
rect 9355 16609 9364 16643
rect 9312 16600 9364 16609
rect 9864 16711 9916 16720
rect 9864 16677 9873 16711
rect 9873 16677 9907 16711
rect 9907 16677 9916 16711
rect 9864 16668 9916 16677
rect 9680 16600 9732 16652
rect 14832 16643 14884 16652
rect 14832 16609 14841 16643
rect 14841 16609 14875 16643
rect 14875 16609 14884 16643
rect 14832 16600 14884 16609
rect 15476 16668 15528 16720
rect 16212 16668 16264 16720
rect 15016 16643 15068 16652
rect 15016 16609 15025 16643
rect 15025 16609 15059 16643
rect 15059 16609 15068 16643
rect 15016 16600 15068 16609
rect 6460 16507 6512 16516
rect 6460 16473 6469 16507
rect 6469 16473 6503 16507
rect 6503 16473 6512 16507
rect 6460 16464 6512 16473
rect 14464 16464 14516 16516
rect 14924 16464 14976 16516
rect 15384 16600 15436 16652
rect 15844 16532 15896 16584
rect 15936 16575 15988 16584
rect 15936 16541 15945 16575
rect 15945 16541 15979 16575
rect 15979 16541 15988 16575
rect 15936 16532 15988 16541
rect 16120 16600 16172 16652
rect 16672 16600 16724 16652
rect 16764 16600 16816 16652
rect 17316 16668 17368 16720
rect 17132 16643 17184 16652
rect 17132 16609 17141 16643
rect 17141 16609 17175 16643
rect 17175 16609 17184 16643
rect 17132 16600 17184 16609
rect 18420 16643 18472 16652
rect 18420 16609 18429 16643
rect 18429 16609 18463 16643
rect 18463 16609 18472 16643
rect 18420 16600 18472 16609
rect 18604 16643 18656 16652
rect 18604 16609 18613 16643
rect 18613 16609 18647 16643
rect 18647 16609 18656 16643
rect 18604 16600 18656 16609
rect 20076 16668 20128 16720
rect 21272 16779 21324 16788
rect 21272 16745 21281 16779
rect 21281 16745 21315 16779
rect 21315 16745 21324 16779
rect 21272 16736 21324 16745
rect 16580 16464 16632 16516
rect 17316 16532 17368 16584
rect 20536 16600 20588 16652
rect 22744 16668 22796 16720
rect 21732 16643 21784 16652
rect 21732 16609 21741 16643
rect 21741 16609 21775 16643
rect 21775 16609 21784 16643
rect 21732 16600 21784 16609
rect 18328 16464 18380 16516
rect 7196 16396 7248 16448
rect 7748 16396 7800 16448
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 10232 16439 10284 16448
rect 10232 16405 10241 16439
rect 10241 16405 10275 16439
rect 10275 16405 10284 16439
rect 10232 16396 10284 16405
rect 16120 16439 16172 16448
rect 16120 16405 16129 16439
rect 16129 16405 16163 16439
rect 16163 16405 16172 16439
rect 16120 16396 16172 16405
rect 17040 16396 17092 16448
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 5080 16124 5132 16176
rect 7104 16192 7156 16244
rect 7472 16124 7524 16176
rect 6920 16099 6972 16108
rect 6920 16065 6929 16099
rect 6929 16065 6963 16099
rect 6963 16065 6972 16099
rect 6920 16056 6972 16065
rect 7196 16056 7248 16108
rect 9036 16056 9088 16108
rect 5540 15988 5592 16040
rect 6184 15988 6236 16040
rect 6460 16031 6512 16040
rect 6460 15997 6469 16031
rect 6469 15997 6503 16031
rect 6503 15997 6512 16031
rect 6460 15988 6512 15997
rect 7564 15988 7616 16040
rect 8576 16031 8628 16040
rect 8576 15997 8585 16031
rect 8585 15997 8619 16031
rect 8619 15997 8628 16031
rect 8576 15988 8628 15997
rect 9680 15988 9732 16040
rect 10784 16031 10836 16040
rect 10784 15997 10793 16031
rect 10793 15997 10827 16031
rect 10827 15997 10836 16031
rect 10784 15988 10836 15997
rect 12992 16124 13044 16176
rect 4804 15920 4856 15972
rect 5632 15920 5684 15972
rect 8116 15852 8168 15904
rect 10324 15920 10376 15972
rect 12532 16031 12584 16040
rect 12532 15997 12541 16031
rect 12541 15997 12575 16031
rect 12575 15997 12584 16031
rect 12532 15988 12584 15997
rect 12992 16031 13044 16040
rect 12992 15997 13001 16031
rect 13001 15997 13035 16031
rect 13035 15997 13044 16031
rect 12992 15988 13044 15997
rect 12256 15920 12308 15972
rect 14832 16192 14884 16244
rect 15016 16192 15068 16244
rect 15476 16235 15528 16244
rect 15476 16201 15485 16235
rect 15485 16201 15519 16235
rect 15519 16201 15528 16235
rect 15476 16192 15528 16201
rect 16672 16192 16724 16244
rect 16856 16192 16908 16244
rect 17500 16192 17552 16244
rect 19432 16235 19484 16244
rect 19432 16201 19441 16235
rect 19441 16201 19475 16235
rect 19475 16201 19484 16235
rect 19432 16192 19484 16201
rect 20352 16192 20404 16244
rect 14832 16056 14884 16108
rect 14464 15988 14516 16040
rect 11980 15852 12032 15904
rect 12900 15895 12952 15904
rect 12900 15861 12909 15895
rect 12909 15861 12943 15895
rect 12943 15861 12952 15895
rect 12900 15852 12952 15861
rect 14740 15988 14792 16040
rect 15108 16056 15160 16108
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 16212 15988 16264 16040
rect 16488 16031 16540 16040
rect 16488 15997 16497 16031
rect 16497 15997 16531 16031
rect 16531 15997 16540 16031
rect 16488 15988 16540 15997
rect 16948 16031 17000 16040
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 17040 16031 17092 16040
rect 17040 15997 17049 16031
rect 17049 15997 17083 16031
rect 17083 15997 17092 16031
rect 17040 15988 17092 15997
rect 17684 15988 17736 16040
rect 18880 15988 18932 16040
rect 19432 16056 19484 16108
rect 19524 16031 19576 16040
rect 19524 15997 19533 16031
rect 19533 15997 19567 16031
rect 19567 15997 19576 16031
rect 19524 15988 19576 15997
rect 20076 16031 20128 16040
rect 20076 15997 20085 16031
rect 20085 15997 20119 16031
rect 20119 15997 20128 16031
rect 20076 15988 20128 15997
rect 15292 15920 15344 15972
rect 17500 15920 17552 15972
rect 20904 15988 20956 16040
rect 21732 16124 21784 16176
rect 22284 16192 22336 16244
rect 21732 16031 21784 16040
rect 21732 15997 21741 16031
rect 21741 15997 21775 16031
rect 21775 15997 21784 16031
rect 21732 15988 21784 15997
rect 21456 15920 21508 15972
rect 22284 15988 22336 16040
rect 22652 15988 22704 16040
rect 14372 15852 14424 15904
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 16764 15895 16816 15904
rect 16764 15861 16773 15895
rect 16773 15861 16807 15895
rect 16807 15861 16816 15895
rect 16764 15852 16816 15861
rect 19708 15895 19760 15904
rect 19708 15861 19717 15895
rect 19717 15861 19751 15895
rect 19751 15861 19760 15895
rect 19708 15852 19760 15861
rect 19892 15852 19944 15904
rect 20352 15895 20404 15904
rect 20352 15861 20361 15895
rect 20361 15861 20395 15895
rect 20395 15861 20404 15895
rect 20352 15852 20404 15861
rect 20444 15852 20496 15904
rect 22100 15920 22152 15972
rect 22560 15895 22612 15904
rect 22560 15861 22569 15895
rect 22569 15861 22603 15895
rect 22603 15861 22612 15895
rect 22560 15852 22612 15861
rect 22836 15852 22888 15904
rect 4322 15750 4374 15802
rect 4386 15750 4438 15802
rect 4450 15750 4502 15802
rect 4514 15750 4566 15802
rect 4578 15750 4630 15802
rect 4896 15580 4948 15632
rect 7564 15691 7616 15700
rect 7564 15657 7573 15691
rect 7573 15657 7607 15691
rect 7607 15657 7616 15691
rect 7564 15648 7616 15657
rect 10416 15648 10468 15700
rect 7748 15623 7800 15632
rect 7748 15589 7757 15623
rect 7757 15589 7791 15623
rect 7791 15589 7800 15623
rect 7748 15580 7800 15589
rect 5080 15555 5132 15564
rect 5080 15521 5089 15555
rect 5089 15521 5123 15555
rect 5123 15521 5132 15555
rect 5080 15512 5132 15521
rect 5632 15512 5684 15564
rect 6368 15512 6420 15564
rect 7472 15555 7524 15564
rect 7472 15521 7481 15555
rect 7481 15521 7515 15555
rect 7515 15521 7524 15555
rect 7472 15512 7524 15521
rect 5816 15487 5868 15496
rect 5816 15453 5825 15487
rect 5825 15453 5859 15487
rect 5859 15453 5868 15487
rect 5816 15444 5868 15453
rect 8116 15555 8168 15564
rect 8116 15521 8125 15555
rect 8125 15521 8159 15555
rect 8159 15521 8168 15555
rect 8116 15512 8168 15521
rect 9036 15512 9088 15564
rect 9680 15555 9732 15564
rect 9680 15521 9690 15555
rect 9690 15521 9724 15555
rect 9724 15521 9732 15555
rect 9680 15512 9732 15521
rect 10324 15512 10376 15564
rect 10784 15648 10836 15700
rect 12256 15648 12308 15700
rect 11336 15580 11388 15632
rect 11520 15512 11572 15564
rect 11888 15555 11940 15564
rect 11888 15521 11897 15555
rect 11897 15521 11931 15555
rect 11931 15521 11940 15555
rect 11888 15512 11940 15521
rect 11980 15555 12032 15564
rect 11980 15521 11989 15555
rect 11989 15521 12023 15555
rect 12023 15521 12032 15555
rect 11980 15512 12032 15521
rect 10140 15419 10192 15428
rect 10140 15385 10149 15419
rect 10149 15385 10183 15419
rect 10183 15385 10192 15419
rect 10140 15376 10192 15385
rect 10692 15444 10744 15496
rect 12256 15555 12308 15564
rect 12256 15521 12265 15555
rect 12265 15521 12299 15555
rect 12299 15521 12308 15555
rect 12256 15512 12308 15521
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 17500 15691 17552 15700
rect 17500 15657 17509 15691
rect 17509 15657 17543 15691
rect 17543 15657 17552 15691
rect 17500 15648 17552 15657
rect 20444 15648 20496 15700
rect 12716 15512 12768 15564
rect 12900 15512 12952 15564
rect 15292 15580 15344 15632
rect 16672 15580 16724 15632
rect 20904 15580 20956 15632
rect 14740 15555 14792 15564
rect 14740 15521 14749 15555
rect 14749 15521 14783 15555
rect 14783 15521 14792 15555
rect 14740 15512 14792 15521
rect 17408 15512 17460 15564
rect 17684 15555 17736 15564
rect 17684 15521 17693 15555
rect 17693 15521 17727 15555
rect 17727 15521 17736 15555
rect 17684 15512 17736 15521
rect 17868 15555 17920 15564
rect 17868 15521 17877 15555
rect 17877 15521 17911 15555
rect 17911 15521 17920 15555
rect 17868 15512 17920 15521
rect 19524 15512 19576 15564
rect 19708 15555 19760 15564
rect 19708 15521 19717 15555
rect 19717 15521 19751 15555
rect 19751 15521 19760 15555
rect 19708 15512 19760 15521
rect 19892 15555 19944 15564
rect 19892 15521 19901 15555
rect 19901 15521 19935 15555
rect 19935 15521 19944 15555
rect 19892 15512 19944 15521
rect 20536 15555 20588 15564
rect 20536 15521 20545 15555
rect 20545 15521 20579 15555
rect 20579 15521 20588 15555
rect 20536 15512 20588 15521
rect 13820 15487 13872 15496
rect 13820 15453 13829 15487
rect 13829 15453 13863 15487
rect 13863 15453 13872 15487
rect 13820 15444 13872 15453
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 18880 15487 18932 15496
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 20628 15487 20680 15496
rect 20628 15453 20637 15487
rect 20637 15453 20671 15487
rect 20671 15453 20680 15487
rect 20628 15444 20680 15453
rect 11888 15376 11940 15428
rect 21732 15512 21784 15564
rect 22652 15512 22704 15564
rect 21456 15444 21508 15496
rect 22100 15444 22152 15496
rect 22008 15376 22060 15428
rect 6552 15308 6604 15360
rect 11336 15308 11388 15360
rect 11520 15351 11572 15360
rect 11520 15317 11529 15351
rect 11529 15317 11563 15351
rect 11563 15317 11572 15351
rect 11520 15308 11572 15317
rect 11612 15308 11664 15360
rect 13544 15308 13596 15360
rect 17776 15351 17828 15360
rect 17776 15317 17785 15351
rect 17785 15317 17819 15351
rect 17819 15317 17828 15351
rect 17776 15308 17828 15317
rect 18420 15351 18472 15360
rect 18420 15317 18429 15351
rect 18429 15317 18463 15351
rect 18463 15317 18472 15351
rect 18420 15308 18472 15317
rect 19800 15351 19852 15360
rect 19800 15317 19809 15351
rect 19809 15317 19843 15351
rect 19843 15317 19852 15351
rect 19800 15308 19852 15317
rect 20352 15308 20404 15360
rect 20628 15351 20680 15360
rect 20628 15317 20637 15351
rect 20637 15317 20671 15351
rect 20671 15317 20680 15351
rect 20628 15308 20680 15317
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 22376 15308 22428 15360
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 10968 15147 11020 15156
rect 10968 15113 10977 15147
rect 10977 15113 11011 15147
rect 11011 15113 11020 15147
rect 10968 15104 11020 15113
rect 11980 15104 12032 15156
rect 12532 15104 12584 15156
rect 13820 15104 13872 15156
rect 9404 15036 9456 15088
rect 9220 15011 9272 15020
rect 9220 14977 9229 15011
rect 9229 14977 9263 15011
rect 9263 14977 9272 15011
rect 9220 14968 9272 14977
rect 9772 14968 9824 15020
rect 13084 15079 13136 15088
rect 13084 15045 13093 15079
rect 13093 15045 13127 15079
rect 13127 15045 13136 15079
rect 13084 15036 13136 15045
rect 9128 14900 9180 14952
rect 9404 14943 9456 14952
rect 9404 14909 9414 14943
rect 9414 14909 9448 14943
rect 9448 14909 9456 14943
rect 9404 14900 9456 14909
rect 9956 14900 10008 14952
rect 10324 14900 10376 14952
rect 14648 15104 14700 15156
rect 17684 15104 17736 15156
rect 15200 15036 15252 15088
rect 14096 14968 14148 15020
rect 11520 14900 11572 14952
rect 10140 14832 10192 14884
rect 9772 14764 9824 14816
rect 10600 14807 10652 14816
rect 10600 14773 10609 14807
rect 10609 14773 10643 14807
rect 10643 14773 10652 14807
rect 10600 14764 10652 14773
rect 11336 14832 11388 14884
rect 13544 14943 13596 14952
rect 13544 14909 13553 14943
rect 13553 14909 13587 14943
rect 13587 14909 13596 14943
rect 13544 14900 13596 14909
rect 12716 14875 12768 14884
rect 12716 14841 12725 14875
rect 12725 14841 12759 14875
rect 12759 14841 12768 14875
rect 12716 14832 12768 14841
rect 12900 14875 12952 14884
rect 12900 14841 12925 14875
rect 12925 14841 12952 14875
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 12900 14832 12952 14841
rect 10876 14764 10928 14816
rect 11428 14764 11480 14816
rect 11796 14764 11848 14816
rect 11888 14807 11940 14816
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 12348 14807 12400 14816
rect 12348 14773 12357 14807
rect 12357 14773 12391 14807
rect 12391 14773 12400 14807
rect 12348 14764 12400 14773
rect 14648 14764 14700 14816
rect 15476 14900 15528 14952
rect 16120 14900 16172 14952
rect 16764 14943 16816 14952
rect 16764 14909 16798 14943
rect 16798 14909 16816 14943
rect 16764 14900 16816 14909
rect 17868 14832 17920 14884
rect 17592 14764 17644 14816
rect 18880 15104 18932 15156
rect 19248 15104 19300 15156
rect 20628 15104 20680 15156
rect 19800 15011 19852 15020
rect 19800 14977 19809 15011
rect 19809 14977 19843 15011
rect 19843 14977 19852 15011
rect 19800 14968 19852 14977
rect 20720 14968 20772 15020
rect 21272 14968 21324 15020
rect 19892 14943 19944 14952
rect 19892 14909 19901 14943
rect 19901 14909 19935 14943
rect 19935 14909 19944 14943
rect 19892 14900 19944 14909
rect 20444 14943 20496 14952
rect 20444 14909 20453 14943
rect 20453 14909 20487 14943
rect 20487 14909 20496 14943
rect 20444 14900 20496 14909
rect 21456 14943 21508 14952
rect 21456 14909 21465 14943
rect 21465 14909 21499 14943
rect 21499 14909 21508 14943
rect 21456 14900 21508 14909
rect 22008 14943 22060 14952
rect 22008 14909 22017 14943
rect 22017 14909 22051 14943
rect 22051 14909 22060 14943
rect 22008 14900 22060 14909
rect 22376 14943 22428 14952
rect 22376 14909 22385 14943
rect 22385 14909 22419 14943
rect 22419 14909 22428 14943
rect 22376 14900 22428 14909
rect 18696 14875 18748 14884
rect 18696 14841 18705 14875
rect 18705 14841 18739 14875
rect 18739 14841 18748 14875
rect 18696 14832 18748 14841
rect 18880 14875 18932 14884
rect 18880 14841 18889 14875
rect 18889 14841 18923 14875
rect 18923 14841 18932 14875
rect 18880 14832 18932 14841
rect 20352 14832 20404 14884
rect 20904 14832 20956 14884
rect 22560 14832 22612 14884
rect 19064 14807 19116 14816
rect 19064 14773 19073 14807
rect 19073 14773 19107 14807
rect 19107 14773 19116 14807
rect 19064 14764 19116 14773
rect 22468 14807 22520 14816
rect 22468 14773 22477 14807
rect 22477 14773 22511 14807
rect 22511 14773 22520 14807
rect 22468 14764 22520 14773
rect 4322 14662 4374 14714
rect 4386 14662 4438 14714
rect 4450 14662 4502 14714
rect 4514 14662 4566 14714
rect 4578 14662 4630 14714
rect 6184 14603 6236 14612
rect 6184 14569 6193 14603
rect 6193 14569 6227 14603
rect 6227 14569 6236 14603
rect 6184 14560 6236 14569
rect 10140 14560 10192 14612
rect 10968 14560 11020 14612
rect 9680 14535 9732 14544
rect 9680 14501 9689 14535
rect 9689 14501 9723 14535
rect 9723 14501 9732 14535
rect 9680 14492 9732 14501
rect 11888 14560 11940 14612
rect 13176 14560 13228 14612
rect 14372 14560 14424 14612
rect 11336 14535 11388 14544
rect 11336 14501 11345 14535
rect 11345 14501 11379 14535
rect 11379 14501 11388 14535
rect 11336 14492 11388 14501
rect 6460 14424 6512 14476
rect 9220 14467 9272 14476
rect 9220 14433 9229 14467
rect 9229 14433 9263 14467
rect 9263 14433 9272 14467
rect 9220 14424 9272 14433
rect 9404 14467 9456 14476
rect 9404 14433 9413 14467
rect 9413 14433 9447 14467
rect 9447 14433 9456 14467
rect 9404 14424 9456 14433
rect 9588 14424 9640 14476
rect 10048 14424 10100 14476
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 10232 14424 10284 14433
rect 6368 14399 6420 14408
rect 6368 14365 6377 14399
rect 6377 14365 6411 14399
rect 6411 14365 6420 14399
rect 6368 14356 6420 14365
rect 9036 14356 9088 14408
rect 9772 14356 9824 14408
rect 10876 14424 10928 14476
rect 11612 14467 11664 14476
rect 11612 14433 11621 14467
rect 11621 14433 11655 14467
rect 11655 14433 11664 14467
rect 11612 14424 11664 14433
rect 12348 14424 12400 14476
rect 11428 14356 11480 14408
rect 13084 14467 13136 14476
rect 13084 14433 13093 14467
rect 13093 14433 13127 14467
rect 13127 14433 13136 14467
rect 13084 14424 13136 14433
rect 13452 14424 13504 14476
rect 14648 14492 14700 14544
rect 15016 14603 15068 14612
rect 15016 14569 15025 14603
rect 15025 14569 15059 14603
rect 15059 14569 15068 14603
rect 15016 14560 15068 14569
rect 18696 14560 18748 14612
rect 18880 14560 18932 14612
rect 21824 14560 21876 14612
rect 14096 14467 14148 14476
rect 14096 14433 14105 14467
rect 14105 14433 14139 14467
rect 14139 14433 14148 14467
rect 14096 14424 14148 14433
rect 17592 14535 17644 14544
rect 17592 14501 17601 14535
rect 17601 14501 17635 14535
rect 17635 14501 17644 14535
rect 17592 14492 17644 14501
rect 16580 14424 16632 14476
rect 17408 14467 17460 14476
rect 17408 14433 17417 14467
rect 17417 14433 17451 14467
rect 17451 14433 17460 14467
rect 17408 14424 17460 14433
rect 17684 14467 17736 14476
rect 17684 14433 17693 14467
rect 17693 14433 17727 14467
rect 17727 14433 17736 14467
rect 17684 14424 17736 14433
rect 10232 14288 10284 14340
rect 12348 14288 12400 14340
rect 16948 14399 17000 14408
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 16948 14356 17000 14365
rect 17500 14356 17552 14408
rect 17960 14467 18012 14476
rect 17960 14433 17969 14467
rect 17969 14433 18003 14467
rect 18003 14433 18012 14467
rect 17960 14424 18012 14433
rect 18604 14467 18656 14476
rect 18604 14433 18613 14467
rect 18613 14433 18647 14467
rect 18647 14433 18656 14467
rect 18604 14424 18656 14433
rect 18052 14356 18104 14408
rect 18144 14399 18196 14408
rect 18144 14365 18153 14399
rect 18153 14365 18187 14399
rect 18187 14365 18196 14399
rect 18144 14356 18196 14365
rect 18420 14356 18472 14408
rect 22100 14492 22152 14544
rect 22928 14492 22980 14544
rect 21548 14467 21600 14476
rect 21548 14433 21557 14467
rect 21557 14433 21591 14467
rect 21591 14433 21600 14467
rect 21548 14424 21600 14433
rect 22376 14424 22428 14476
rect 22744 14467 22796 14476
rect 22744 14433 22779 14467
rect 22779 14433 22796 14467
rect 22744 14424 22796 14433
rect 6000 14220 6052 14272
rect 9956 14220 10008 14272
rect 10140 14263 10192 14272
rect 10140 14229 10149 14263
rect 10149 14229 10183 14263
rect 10183 14229 10192 14263
rect 10140 14220 10192 14229
rect 10876 14220 10928 14272
rect 11796 14263 11848 14272
rect 11796 14229 11805 14263
rect 11805 14229 11839 14263
rect 11839 14229 11848 14263
rect 11796 14220 11848 14229
rect 13728 14220 13780 14272
rect 14280 14263 14332 14272
rect 14280 14229 14289 14263
rect 14289 14229 14323 14263
rect 14323 14229 14332 14263
rect 14280 14220 14332 14229
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 18328 14288 18380 14340
rect 14648 14220 14700 14272
rect 16764 14263 16816 14272
rect 16764 14229 16773 14263
rect 16773 14229 16807 14263
rect 16807 14229 16816 14263
rect 16764 14220 16816 14229
rect 17408 14220 17460 14272
rect 21916 14399 21968 14408
rect 21916 14365 21925 14399
rect 21925 14365 21959 14399
rect 21959 14365 21968 14399
rect 21916 14356 21968 14365
rect 18972 14220 19024 14272
rect 19248 14263 19300 14272
rect 19248 14229 19257 14263
rect 19257 14229 19291 14263
rect 19291 14229 19300 14263
rect 19248 14220 19300 14229
rect 19340 14220 19392 14272
rect 20812 14220 20864 14272
rect 22468 14288 22520 14340
rect 22836 14288 22888 14340
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 6184 14016 6236 14068
rect 9588 14016 9640 14068
rect 5540 13812 5592 13864
rect 9220 13948 9272 14000
rect 10048 13948 10100 14000
rect 7656 13923 7708 13932
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 8116 13880 8168 13932
rect 7104 13855 7156 13864
rect 7104 13821 7113 13855
rect 7113 13821 7147 13855
rect 7147 13821 7156 13855
rect 7104 13812 7156 13821
rect 7012 13744 7064 13796
rect 5816 13676 5868 13728
rect 7104 13676 7156 13728
rect 9036 13812 9088 13864
rect 9404 13812 9456 13864
rect 9772 13855 9824 13864
rect 9772 13821 9781 13855
rect 9781 13821 9815 13855
rect 9815 13821 9824 13855
rect 9772 13812 9824 13821
rect 9956 13855 10008 13864
rect 9956 13821 9965 13855
rect 9965 13821 9999 13855
rect 9999 13821 10008 13855
rect 9956 13812 10008 13821
rect 10600 13855 10652 13864
rect 10600 13821 10609 13855
rect 10609 13821 10643 13855
rect 10643 13821 10652 13855
rect 10600 13812 10652 13821
rect 11336 14016 11388 14068
rect 14648 14059 14700 14068
rect 14648 14025 14657 14059
rect 14657 14025 14691 14059
rect 14691 14025 14700 14059
rect 14648 14016 14700 14025
rect 16948 14059 17000 14068
rect 16948 14025 16957 14059
rect 16957 14025 16991 14059
rect 16991 14025 17000 14059
rect 16948 14016 17000 14025
rect 17868 14016 17920 14068
rect 17960 14059 18012 14068
rect 17960 14025 17969 14059
rect 17969 14025 18003 14059
rect 18003 14025 18012 14059
rect 17960 14016 18012 14025
rect 18052 14059 18104 14068
rect 18052 14025 18061 14059
rect 18061 14025 18095 14059
rect 18095 14025 18104 14059
rect 18052 14016 18104 14025
rect 19064 14059 19116 14068
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 20536 14016 20588 14068
rect 21456 14016 21508 14068
rect 21916 14059 21968 14068
rect 21916 14025 21925 14059
rect 21925 14025 21959 14059
rect 21959 14025 21968 14059
rect 21916 14016 21968 14025
rect 13820 13948 13872 14000
rect 12348 13880 12400 13932
rect 13176 13923 13228 13932
rect 13176 13889 13185 13923
rect 13185 13889 13219 13923
rect 13219 13889 13228 13923
rect 13176 13880 13228 13889
rect 13268 13923 13320 13932
rect 13268 13889 13277 13923
rect 13277 13889 13311 13923
rect 13311 13889 13320 13923
rect 13268 13880 13320 13889
rect 10968 13812 11020 13864
rect 12992 13855 13044 13864
rect 12992 13821 13001 13855
rect 13001 13821 13035 13855
rect 13035 13821 13044 13855
rect 12992 13812 13044 13821
rect 13728 13855 13780 13864
rect 13728 13821 13737 13855
rect 13737 13821 13771 13855
rect 13771 13821 13780 13855
rect 13728 13812 13780 13821
rect 14096 13812 14148 13864
rect 14372 13812 14424 13864
rect 14924 13880 14976 13932
rect 15476 13855 15528 13864
rect 15476 13821 15485 13855
rect 15485 13821 15519 13855
rect 15519 13821 15528 13855
rect 15476 13812 15528 13821
rect 19340 13948 19392 14000
rect 18144 13880 18196 13932
rect 19984 13880 20036 13932
rect 16764 13812 16816 13864
rect 13084 13744 13136 13796
rect 16120 13744 16172 13796
rect 18328 13855 18380 13864
rect 9496 13676 9548 13728
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 10416 13719 10468 13728
rect 10416 13685 10425 13719
rect 10425 13685 10459 13719
rect 10459 13685 10468 13719
rect 10416 13676 10468 13685
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 14096 13719 14148 13728
rect 14096 13685 14105 13719
rect 14105 13685 14139 13719
rect 14139 13685 14148 13719
rect 14096 13676 14148 13685
rect 16580 13676 16632 13728
rect 17592 13787 17644 13796
rect 17592 13753 17601 13787
rect 17601 13753 17635 13787
rect 17635 13753 17644 13787
rect 17592 13744 17644 13753
rect 18328 13821 18337 13855
rect 18337 13821 18371 13855
rect 18371 13821 18380 13855
rect 18328 13812 18380 13821
rect 18788 13855 18840 13864
rect 18788 13821 18797 13855
rect 18797 13821 18831 13855
rect 18831 13821 18840 13855
rect 18788 13812 18840 13821
rect 18972 13812 19024 13864
rect 19892 13812 19944 13864
rect 17960 13676 18012 13728
rect 19892 13719 19944 13728
rect 19892 13685 19901 13719
rect 19901 13685 19935 13719
rect 19935 13685 19944 13719
rect 19892 13676 19944 13685
rect 20260 13855 20312 13864
rect 20260 13821 20269 13855
rect 20269 13821 20303 13855
rect 20303 13821 20312 13855
rect 20260 13812 20312 13821
rect 21088 13812 21140 13864
rect 22100 13855 22152 13864
rect 22100 13821 22109 13855
rect 22109 13821 22143 13855
rect 22143 13821 22152 13855
rect 22100 13812 22152 13821
rect 22284 13812 22336 13864
rect 20536 13676 20588 13728
rect 22100 13676 22152 13728
rect 4322 13574 4374 13626
rect 4386 13574 4438 13626
rect 4450 13574 4502 13626
rect 4514 13574 4566 13626
rect 4578 13574 4630 13626
rect 5540 13472 5592 13524
rect 6184 13515 6236 13524
rect 6184 13481 6193 13515
rect 6193 13481 6227 13515
rect 6227 13481 6236 13515
rect 6184 13472 6236 13481
rect 5724 13404 5776 13456
rect 8116 13404 8168 13456
rect 7104 13336 7156 13388
rect 7288 13379 7340 13388
rect 7288 13345 7322 13379
rect 7322 13345 7340 13379
rect 7288 13336 7340 13345
rect 10140 13472 10192 13524
rect 9496 13404 9548 13456
rect 9220 13379 9272 13388
rect 9220 13345 9229 13379
rect 9229 13345 9263 13379
rect 9263 13345 9272 13379
rect 9220 13336 9272 13345
rect 9312 13379 9364 13388
rect 9312 13345 9321 13379
rect 9321 13345 9355 13379
rect 9355 13345 9364 13379
rect 9312 13336 9364 13345
rect 9588 13379 9640 13388
rect 9588 13345 9597 13379
rect 9597 13345 9631 13379
rect 9631 13345 9640 13379
rect 9588 13336 9640 13345
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 11796 13379 11848 13388
rect 11796 13345 11805 13379
rect 11805 13345 11839 13379
rect 11839 13345 11848 13379
rect 11796 13336 11848 13345
rect 12348 13472 12400 13524
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 13268 13472 13320 13524
rect 16120 13515 16172 13524
rect 16120 13481 16129 13515
rect 16129 13481 16163 13515
rect 16163 13481 16172 13515
rect 16120 13472 16172 13481
rect 18144 13472 18196 13524
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 12072 13311 12124 13320
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 12808 13379 12860 13388
rect 12808 13345 12817 13379
rect 12817 13345 12851 13379
rect 12851 13345 12860 13379
rect 12808 13336 12860 13345
rect 13728 13336 13780 13388
rect 14096 13336 14148 13388
rect 14372 13379 14424 13388
rect 14372 13345 14381 13379
rect 14381 13345 14415 13379
rect 14415 13345 14424 13379
rect 14372 13336 14424 13345
rect 12532 13268 12584 13320
rect 13912 13268 13964 13320
rect 14832 13336 14884 13388
rect 16580 13404 16632 13456
rect 17408 13404 17460 13456
rect 17868 13404 17920 13456
rect 19248 13404 19300 13456
rect 20720 13404 20772 13456
rect 20904 13404 20956 13456
rect 21180 13404 21232 13456
rect 9312 13200 9364 13252
rect 20168 13336 20220 13388
rect 21640 13336 21692 13388
rect 22100 13404 22152 13456
rect 22928 13404 22980 13456
rect 15292 13268 15344 13320
rect 16396 13268 16448 13320
rect 16856 13268 16908 13320
rect 16488 13200 16540 13252
rect 19340 13200 19392 13252
rect 20536 13311 20588 13320
rect 20536 13277 20545 13311
rect 20545 13277 20579 13311
rect 20579 13277 20588 13311
rect 20536 13268 20588 13277
rect 20628 13311 20680 13320
rect 20628 13277 20637 13311
rect 20637 13277 20671 13311
rect 20671 13277 20680 13311
rect 20628 13268 20680 13277
rect 20812 13268 20864 13320
rect 21824 13268 21876 13320
rect 22192 13311 22244 13320
rect 22192 13277 22201 13311
rect 22201 13277 22235 13311
rect 22235 13277 22244 13311
rect 22192 13268 22244 13277
rect 8392 13175 8444 13184
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 9036 13175 9088 13184
rect 9036 13141 9045 13175
rect 9045 13141 9079 13175
rect 9079 13141 9088 13175
rect 9036 13132 9088 13141
rect 10140 13175 10192 13184
rect 10140 13141 10149 13175
rect 10149 13141 10183 13175
rect 10183 13141 10192 13175
rect 10140 13132 10192 13141
rect 11612 13175 11664 13184
rect 11612 13141 11621 13175
rect 11621 13141 11655 13175
rect 11655 13141 11664 13175
rect 11612 13132 11664 13141
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 14188 13132 14240 13184
rect 18604 13132 18656 13184
rect 19708 13175 19760 13184
rect 19708 13141 19717 13175
rect 19717 13141 19751 13175
rect 19751 13141 19760 13175
rect 19708 13132 19760 13141
rect 19892 13175 19944 13184
rect 19892 13141 19901 13175
rect 19901 13141 19935 13175
rect 19935 13141 19944 13175
rect 19892 13132 19944 13141
rect 20260 13132 20312 13184
rect 20812 13132 20864 13184
rect 21272 13132 21324 13184
rect 21456 13175 21508 13184
rect 21456 13141 21465 13175
rect 21465 13141 21499 13175
rect 21499 13141 21508 13175
rect 21456 13132 21508 13141
rect 21640 13175 21692 13184
rect 21640 13141 21649 13175
rect 21649 13141 21683 13175
rect 21683 13141 21692 13175
rect 21640 13132 21692 13141
rect 22376 13200 22428 13252
rect 22652 13243 22704 13252
rect 22652 13209 22661 13243
rect 22661 13209 22695 13243
rect 22695 13209 22704 13243
rect 22652 13200 22704 13209
rect 22100 13175 22152 13184
rect 22100 13141 22109 13175
rect 22109 13141 22143 13175
rect 22143 13141 22152 13175
rect 22100 13132 22152 13141
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 6368 12928 6420 12980
rect 6552 12971 6604 12980
rect 6552 12937 6561 12971
rect 6561 12937 6595 12971
rect 6595 12937 6604 12971
rect 6552 12928 6604 12937
rect 7288 12928 7340 12980
rect 7104 12860 7156 12912
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 11060 12928 11112 12980
rect 12072 12928 12124 12980
rect 15292 12971 15344 12980
rect 15292 12937 15301 12971
rect 15301 12937 15335 12971
rect 15335 12937 15344 12971
rect 15292 12928 15344 12937
rect 20536 12928 20588 12980
rect 20996 12971 21048 12980
rect 20996 12937 21005 12971
rect 21005 12937 21039 12971
rect 21039 12937 21048 12971
rect 20996 12928 21048 12937
rect 21088 12971 21140 12980
rect 21088 12937 21097 12971
rect 21097 12937 21131 12971
rect 21131 12937 21140 12971
rect 21088 12928 21140 12937
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 14924 12860 14976 12912
rect 8116 12792 8168 12801
rect 10140 12792 10192 12844
rect 6000 12767 6052 12776
rect 6000 12733 6018 12767
rect 6018 12733 6052 12767
rect 6000 12724 6052 12733
rect 6184 12656 6236 12708
rect 6552 12767 6604 12776
rect 6552 12733 6561 12767
rect 6561 12733 6595 12767
rect 6595 12733 6604 12767
rect 6552 12724 6604 12733
rect 8392 12724 8444 12776
rect 8668 12724 8720 12776
rect 10416 12767 10468 12776
rect 10416 12733 10425 12767
rect 10425 12733 10459 12767
rect 10459 12733 10468 12767
rect 10416 12724 10468 12733
rect 8484 12656 8536 12708
rect 9036 12656 9088 12708
rect 9220 12656 9272 12708
rect 15568 12792 15620 12844
rect 19340 12860 19392 12912
rect 22192 12860 22244 12912
rect 16856 12792 16908 12844
rect 12348 12724 12400 12776
rect 12716 12724 12768 12776
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 14188 12767 14240 12776
rect 14188 12733 14222 12767
rect 14222 12733 14240 12767
rect 12624 12656 12676 12708
rect 14188 12724 14240 12733
rect 18144 12792 18196 12844
rect 17868 12767 17920 12776
rect 17868 12733 17877 12767
rect 17877 12733 17911 12767
rect 17911 12733 17920 12767
rect 17868 12724 17920 12733
rect 15476 12656 15528 12708
rect 18052 12656 18104 12708
rect 18604 12724 18656 12776
rect 19064 12699 19116 12708
rect 19064 12665 19073 12699
rect 19073 12665 19107 12699
rect 19107 12665 19116 12699
rect 19064 12656 19116 12665
rect 19248 12699 19300 12708
rect 19248 12665 19257 12699
rect 19257 12665 19291 12699
rect 19291 12665 19300 12699
rect 19248 12656 19300 12665
rect 5540 12588 5592 12640
rect 7104 12588 7156 12640
rect 8944 12588 8996 12640
rect 9404 12588 9456 12640
rect 11704 12588 11756 12640
rect 12532 12588 12584 12640
rect 12716 12588 12768 12640
rect 15384 12631 15436 12640
rect 15384 12597 15393 12631
rect 15393 12597 15427 12631
rect 15427 12597 15436 12631
rect 15384 12588 15436 12597
rect 15752 12631 15804 12640
rect 15752 12597 15761 12631
rect 15761 12597 15795 12631
rect 15795 12597 15804 12631
rect 15752 12588 15804 12597
rect 17960 12631 18012 12640
rect 17960 12597 17969 12631
rect 17969 12597 18003 12631
rect 18003 12597 18012 12631
rect 17960 12588 18012 12597
rect 18420 12588 18472 12640
rect 19156 12588 19208 12640
rect 19708 12724 19760 12776
rect 21364 12724 21416 12776
rect 21640 12767 21692 12776
rect 21640 12733 21649 12767
rect 21649 12733 21683 12767
rect 21683 12733 21692 12767
rect 21640 12724 21692 12733
rect 19432 12699 19484 12708
rect 19432 12665 19441 12699
rect 19441 12665 19475 12699
rect 19475 12665 19484 12699
rect 19432 12656 19484 12665
rect 21456 12656 21508 12708
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 23020 12767 23072 12776
rect 23020 12733 23029 12767
rect 23029 12733 23063 12767
rect 23063 12733 23072 12767
rect 23020 12724 23072 12733
rect 22928 12656 22980 12708
rect 21732 12631 21784 12640
rect 21732 12597 21741 12631
rect 21741 12597 21775 12631
rect 21775 12597 21784 12631
rect 21732 12588 21784 12597
rect 21916 12631 21968 12640
rect 21916 12597 21925 12631
rect 21925 12597 21959 12631
rect 21959 12597 21968 12631
rect 21916 12588 21968 12597
rect 4322 12486 4374 12538
rect 4386 12486 4438 12538
rect 4450 12486 4502 12538
rect 4514 12486 4566 12538
rect 4578 12486 4630 12538
rect 7196 12384 7248 12436
rect 11152 12384 11204 12436
rect 11980 12384 12032 12436
rect 12624 12384 12676 12436
rect 5540 12316 5592 12368
rect 5724 12316 5776 12368
rect 7012 12316 7064 12368
rect 11612 12359 11664 12368
rect 6736 12291 6788 12300
rect 6736 12257 6745 12291
rect 6745 12257 6779 12291
rect 6779 12257 6788 12291
rect 6736 12248 6788 12257
rect 7104 12291 7156 12300
rect 7104 12257 7113 12291
rect 7113 12257 7147 12291
rect 7147 12257 7156 12291
rect 7104 12248 7156 12257
rect 11612 12325 11646 12359
rect 11646 12325 11664 12359
rect 11612 12316 11664 12325
rect 10232 12248 10284 12300
rect 13360 12248 13412 12300
rect 13820 12248 13872 12300
rect 13912 12291 13964 12300
rect 13912 12257 13921 12291
rect 13921 12257 13955 12291
rect 13955 12257 13964 12291
rect 13912 12248 13964 12257
rect 16580 12316 16632 12368
rect 17868 12384 17920 12436
rect 18604 12384 18656 12436
rect 20720 12384 20772 12436
rect 17960 12359 18012 12368
rect 17960 12325 17994 12359
rect 17994 12325 18012 12359
rect 17960 12316 18012 12325
rect 18144 12316 18196 12368
rect 21732 12316 21784 12368
rect 18236 12248 18288 12300
rect 20812 12291 20864 12300
rect 20812 12257 20821 12291
rect 20821 12257 20855 12291
rect 20855 12257 20864 12291
rect 20812 12248 20864 12257
rect 20996 12291 21048 12300
rect 20996 12257 21005 12291
rect 21005 12257 21039 12291
rect 21039 12257 21048 12291
rect 20996 12248 21048 12257
rect 21088 12248 21140 12300
rect 22652 12248 22704 12300
rect 6368 12180 6420 12232
rect 6184 12112 6236 12164
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 11336 12223 11388 12232
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11336 12180 11388 12189
rect 7472 12112 7524 12164
rect 5816 12087 5868 12096
rect 5816 12053 5825 12087
rect 5825 12053 5859 12087
rect 5859 12053 5868 12087
rect 5816 12044 5868 12053
rect 6368 12044 6420 12096
rect 7380 12044 7432 12096
rect 9864 12044 9916 12096
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 16580 12223 16632 12232
rect 16580 12189 16589 12223
rect 16589 12189 16623 12223
rect 16623 12189 16632 12223
rect 16580 12180 16632 12189
rect 16764 12180 16816 12232
rect 15108 12112 15160 12164
rect 19156 12223 19208 12232
rect 19156 12189 19165 12223
rect 19165 12189 19199 12223
rect 19199 12189 19208 12223
rect 19156 12180 19208 12189
rect 21272 12180 21324 12232
rect 14832 12044 14884 12096
rect 16120 12044 16172 12096
rect 16856 12087 16908 12096
rect 16856 12053 16865 12087
rect 16865 12053 16899 12087
rect 16899 12053 16908 12087
rect 16856 12044 16908 12053
rect 17960 12044 18012 12096
rect 19064 12044 19116 12096
rect 21456 12087 21508 12096
rect 21456 12053 21465 12087
rect 21465 12053 21499 12087
rect 21499 12053 21508 12087
rect 21456 12044 21508 12053
rect 21640 12044 21692 12096
rect 21916 12044 21968 12096
rect 22928 12044 22980 12096
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 7104 11840 7156 11892
rect 15752 11840 15804 11892
rect 6920 11815 6972 11824
rect 6920 11781 6929 11815
rect 6929 11781 6963 11815
rect 6963 11781 6972 11815
rect 6920 11772 6972 11781
rect 5816 11704 5868 11756
rect 6644 11704 6696 11756
rect 7472 11704 7524 11756
rect 8300 11704 8352 11756
rect 6000 11679 6052 11688
rect 6000 11645 6009 11679
rect 6009 11645 6043 11679
rect 6043 11645 6052 11679
rect 6000 11636 6052 11645
rect 6460 11611 6512 11620
rect 6460 11577 6469 11611
rect 6469 11577 6503 11611
rect 6503 11577 6512 11611
rect 6460 11568 6512 11577
rect 7104 11679 7156 11688
rect 7104 11645 7113 11679
rect 7113 11645 7147 11679
rect 7147 11645 7156 11679
rect 7104 11636 7156 11645
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 8392 11636 8444 11688
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 16120 11883 16172 11892
rect 16120 11849 16129 11883
rect 16129 11849 16163 11883
rect 16163 11849 16172 11883
rect 16120 11840 16172 11849
rect 16580 11883 16632 11892
rect 16580 11849 16589 11883
rect 16589 11849 16623 11883
rect 16623 11849 16632 11883
rect 16580 11840 16632 11849
rect 16764 11840 16816 11892
rect 18052 11883 18104 11892
rect 18052 11849 18061 11883
rect 18061 11849 18095 11883
rect 18095 11849 18104 11883
rect 18052 11840 18104 11849
rect 18236 11883 18288 11892
rect 18236 11849 18245 11883
rect 18245 11849 18279 11883
rect 18279 11849 18288 11883
rect 18236 11840 18288 11849
rect 20352 11840 20404 11892
rect 21180 11840 21232 11892
rect 22284 11840 22336 11892
rect 18788 11772 18840 11824
rect 8668 11636 8720 11688
rect 10232 11636 10284 11688
rect 14096 11636 14148 11688
rect 9404 11568 9456 11620
rect 11244 11611 11296 11620
rect 11244 11577 11278 11611
rect 11278 11577 11296 11611
rect 11244 11568 11296 11577
rect 11336 11568 11388 11620
rect 15384 11636 15436 11688
rect 15016 11568 15068 11620
rect 15200 11568 15252 11620
rect 17224 11679 17276 11688
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 17408 11636 17460 11688
rect 6552 11500 6604 11552
rect 6644 11543 6696 11552
rect 6644 11509 6669 11543
rect 6669 11509 6696 11543
rect 6644 11500 6696 11509
rect 6828 11543 6880 11552
rect 6828 11509 6837 11543
rect 6837 11509 6871 11543
rect 6871 11509 6880 11543
rect 6828 11500 6880 11509
rect 7656 11500 7708 11552
rect 8576 11500 8628 11552
rect 9220 11500 9272 11552
rect 10324 11500 10376 11552
rect 12348 11543 12400 11552
rect 12348 11509 12357 11543
rect 12357 11509 12391 11543
rect 12391 11509 12400 11543
rect 12348 11500 12400 11509
rect 15292 11500 15344 11552
rect 16672 11568 16724 11620
rect 19432 11636 19484 11688
rect 21364 11679 21416 11688
rect 21364 11645 21373 11679
rect 21373 11645 21407 11679
rect 21407 11645 21416 11679
rect 21364 11636 21416 11645
rect 17316 11500 17368 11552
rect 17960 11568 18012 11620
rect 18420 11568 18472 11620
rect 19340 11568 19392 11620
rect 19432 11543 19484 11552
rect 21272 11568 21324 11620
rect 22928 11636 22980 11688
rect 21548 11568 21600 11620
rect 19432 11509 19457 11543
rect 19457 11509 19484 11543
rect 19432 11500 19484 11509
rect 22376 11500 22428 11552
rect 4322 11398 4374 11450
rect 4386 11398 4438 11450
rect 4450 11398 4502 11450
rect 4514 11398 4566 11450
rect 4578 11398 4630 11450
rect 7472 11339 7524 11348
rect 7472 11305 7481 11339
rect 7481 11305 7515 11339
rect 7515 11305 7524 11339
rect 7472 11296 7524 11305
rect 9312 11296 9364 11348
rect 9404 11339 9456 11348
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 9864 11339 9916 11348
rect 9864 11305 9873 11339
rect 9873 11305 9907 11339
rect 9907 11305 9916 11339
rect 9864 11296 9916 11305
rect 5632 11228 5684 11280
rect 4620 11092 4672 11144
rect 5724 11160 5776 11212
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 6184 11271 6236 11280
rect 6184 11237 6193 11271
rect 6193 11237 6227 11271
rect 6227 11237 6236 11271
rect 6184 11228 6236 11237
rect 5080 11092 5132 11144
rect 6184 11092 6236 11144
rect 6736 11228 6788 11280
rect 6552 11160 6604 11212
rect 6828 11203 6880 11212
rect 6828 11169 6837 11203
rect 6837 11169 6871 11203
rect 6871 11169 6880 11203
rect 6828 11160 6880 11169
rect 7104 11203 7156 11212
rect 7104 11169 7113 11203
rect 7113 11169 7147 11203
rect 7147 11169 7156 11203
rect 7104 11160 7156 11169
rect 8576 11271 8628 11280
rect 8576 11237 8585 11271
rect 8585 11237 8619 11271
rect 8619 11237 8628 11271
rect 8576 11228 8628 11237
rect 7380 11203 7432 11212
rect 7380 11169 7389 11203
rect 7389 11169 7423 11203
rect 7423 11169 7432 11203
rect 7380 11160 7432 11169
rect 7656 11203 7708 11212
rect 7656 11169 7665 11203
rect 7665 11169 7699 11203
rect 7699 11169 7708 11203
rect 7656 11160 7708 11169
rect 8300 11092 8352 11144
rect 8392 11092 8444 11144
rect 10232 11203 10284 11212
rect 10232 11169 10241 11203
rect 10241 11169 10275 11203
rect 10275 11169 10284 11203
rect 10232 11160 10284 11169
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 11704 11339 11756 11348
rect 11704 11305 11713 11339
rect 11713 11305 11747 11339
rect 11747 11305 11756 11339
rect 11704 11296 11756 11305
rect 10324 11135 10376 11144
rect 8760 11024 8812 11076
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 6920 10956 6972 11008
rect 8300 10956 8352 11008
rect 9496 10956 9548 11008
rect 11152 10956 11204 11008
rect 12532 11203 12584 11212
rect 12532 11169 12541 11203
rect 12541 11169 12575 11203
rect 12575 11169 12584 11203
rect 12532 11160 12584 11169
rect 12716 11203 12768 11212
rect 12716 11169 12725 11203
rect 12725 11169 12759 11203
rect 12759 11169 12768 11203
rect 12716 11160 12768 11169
rect 12348 11092 12400 11144
rect 13728 11160 13780 11212
rect 15200 11160 15252 11212
rect 15292 11203 15344 11212
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 15568 11160 15620 11212
rect 16764 11339 16816 11348
rect 16764 11305 16773 11339
rect 16773 11305 16807 11339
rect 16807 11305 16816 11339
rect 16764 11296 16816 11305
rect 17408 11339 17460 11348
rect 17408 11305 17417 11339
rect 17417 11305 17451 11339
rect 17451 11305 17460 11339
rect 17408 11296 17460 11305
rect 17592 11296 17644 11348
rect 18144 11296 18196 11348
rect 16396 11271 16448 11280
rect 16396 11237 16405 11271
rect 16405 11237 16439 11271
rect 16439 11237 16448 11271
rect 16396 11228 16448 11237
rect 18420 11228 18472 11280
rect 17040 11203 17092 11212
rect 17040 11169 17049 11203
rect 17049 11169 17083 11203
rect 17083 11169 17092 11203
rect 17040 11160 17092 11169
rect 17868 11203 17920 11212
rect 17868 11169 17877 11203
rect 17877 11169 17911 11203
rect 17911 11169 17920 11203
rect 17868 11160 17920 11169
rect 19432 11296 19484 11348
rect 20352 11296 20404 11348
rect 21548 11339 21600 11348
rect 21548 11305 21557 11339
rect 21557 11305 21591 11339
rect 21591 11305 21600 11339
rect 21548 11296 21600 11305
rect 21640 11296 21692 11348
rect 22284 11228 22336 11280
rect 16580 11092 16632 11144
rect 16856 11092 16908 11144
rect 20720 11203 20772 11212
rect 20720 11169 20729 11203
rect 20729 11169 20763 11203
rect 20763 11169 20772 11203
rect 20720 11160 20772 11169
rect 22100 11203 22152 11212
rect 22100 11169 22109 11203
rect 22109 11169 22143 11203
rect 22143 11169 22152 11203
rect 22100 11160 22152 11169
rect 22376 11203 22428 11212
rect 22376 11169 22385 11203
rect 22385 11169 22419 11203
rect 22419 11169 22428 11203
rect 22376 11160 22428 11169
rect 21180 11092 21232 11144
rect 13728 11024 13780 11076
rect 14832 11024 14884 11076
rect 17224 11024 17276 11076
rect 11520 10956 11572 11008
rect 12624 10999 12676 11008
rect 12624 10965 12633 10999
rect 12633 10965 12667 10999
rect 12667 10965 12676 10999
rect 12624 10956 12676 10965
rect 14556 10956 14608 11008
rect 14924 10999 14976 11008
rect 14924 10965 14933 10999
rect 14933 10965 14967 10999
rect 14967 10965 14976 10999
rect 14924 10956 14976 10965
rect 16580 10999 16632 11008
rect 16580 10965 16589 10999
rect 16589 10965 16623 10999
rect 16623 10965 16632 10999
rect 16580 10956 16632 10965
rect 18236 10956 18288 11008
rect 18328 10999 18380 11008
rect 18328 10965 18337 10999
rect 18337 10965 18371 10999
rect 18371 10965 18380 10999
rect 18328 10956 18380 10965
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 6184 10752 6236 10804
rect 7104 10752 7156 10804
rect 9496 10795 9548 10804
rect 9496 10761 9505 10795
rect 9505 10761 9539 10795
rect 9539 10761 9548 10795
rect 9496 10752 9548 10761
rect 3976 10548 4028 10600
rect 4620 10591 4672 10600
rect 4620 10557 4629 10591
rect 4629 10557 4663 10591
rect 4663 10557 4672 10591
rect 4620 10548 4672 10557
rect 4252 10480 4304 10532
rect 4896 10591 4948 10600
rect 4896 10557 4905 10591
rect 4905 10557 4939 10591
rect 4939 10557 4948 10591
rect 4896 10548 4948 10557
rect 8300 10616 8352 10668
rect 8852 10616 8904 10668
rect 9956 10752 10008 10804
rect 10508 10752 10560 10804
rect 12532 10795 12584 10804
rect 12532 10761 12541 10795
rect 12541 10761 12575 10795
rect 12575 10761 12584 10795
rect 12532 10752 12584 10761
rect 18328 10752 18380 10804
rect 20720 10752 20772 10804
rect 22008 10752 22060 10804
rect 10416 10727 10468 10736
rect 10416 10693 10425 10727
rect 10425 10693 10459 10727
rect 10459 10693 10468 10727
rect 10416 10684 10468 10693
rect 5632 10548 5684 10600
rect 6460 10548 6512 10600
rect 8392 10548 8444 10600
rect 5172 10523 5224 10532
rect 5172 10489 5206 10523
rect 5206 10489 5224 10523
rect 5172 10480 5224 10489
rect 6368 10523 6420 10532
rect 6368 10489 6377 10523
rect 6377 10489 6411 10523
rect 6411 10489 6420 10523
rect 6368 10480 6420 10489
rect 9772 10548 9824 10600
rect 10324 10548 10376 10600
rect 10508 10548 10560 10600
rect 4712 10455 4764 10464
rect 4712 10421 4721 10455
rect 4721 10421 4755 10455
rect 4755 10421 4764 10455
rect 4712 10412 4764 10421
rect 6736 10455 6788 10464
rect 6736 10421 6745 10455
rect 6745 10421 6779 10455
rect 6779 10421 6788 10455
rect 6736 10412 6788 10421
rect 9220 10412 9272 10464
rect 9680 10455 9732 10464
rect 9680 10421 9689 10455
rect 9689 10421 9723 10455
rect 9723 10421 9732 10455
rect 9680 10412 9732 10421
rect 10324 10455 10376 10464
rect 10324 10421 10333 10455
rect 10333 10421 10367 10455
rect 10367 10421 10376 10455
rect 10324 10412 10376 10421
rect 11060 10548 11112 10600
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 12624 10684 12676 10736
rect 14556 10659 14608 10668
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 14556 10616 14608 10625
rect 12348 10548 12400 10600
rect 12716 10591 12768 10600
rect 12716 10557 12725 10591
rect 12725 10557 12759 10591
rect 12759 10557 12768 10591
rect 12716 10548 12768 10557
rect 13728 10591 13780 10600
rect 13728 10557 13737 10591
rect 13737 10557 13771 10591
rect 13771 10557 13780 10591
rect 13728 10548 13780 10557
rect 14832 10548 14884 10600
rect 14924 10548 14976 10600
rect 17500 10684 17552 10736
rect 22744 10795 22796 10804
rect 22744 10761 22753 10795
rect 22753 10761 22787 10795
rect 22787 10761 22796 10795
rect 22744 10752 22796 10761
rect 22560 10684 22612 10736
rect 18236 10591 18288 10600
rect 18236 10557 18254 10591
rect 18254 10557 18288 10591
rect 18236 10548 18288 10557
rect 14740 10480 14792 10532
rect 16672 10523 16724 10532
rect 16672 10489 16681 10523
rect 16681 10489 16715 10523
rect 16715 10489 16724 10523
rect 16672 10480 16724 10489
rect 18144 10480 18196 10532
rect 19156 10548 19208 10600
rect 21088 10480 21140 10532
rect 21916 10548 21968 10600
rect 22100 10591 22152 10600
rect 22100 10557 22109 10591
rect 22109 10557 22143 10591
rect 22143 10557 22152 10591
rect 22100 10548 22152 10557
rect 22376 10591 22428 10600
rect 22376 10557 22385 10591
rect 22385 10557 22419 10591
rect 22419 10557 22428 10591
rect 22376 10548 22428 10557
rect 22652 10548 22704 10600
rect 11612 10412 11664 10464
rect 12164 10455 12216 10464
rect 12164 10421 12173 10455
rect 12173 10421 12207 10455
rect 12207 10421 12216 10455
rect 12164 10412 12216 10421
rect 13728 10455 13780 10464
rect 13728 10421 13737 10455
rect 13737 10421 13771 10455
rect 13771 10421 13780 10455
rect 13728 10412 13780 10421
rect 15108 10412 15160 10464
rect 21272 10455 21324 10464
rect 21272 10421 21281 10455
rect 21281 10421 21315 10455
rect 21315 10421 21324 10455
rect 21272 10412 21324 10421
rect 22468 10412 22520 10464
rect 4322 10310 4374 10362
rect 4386 10310 4438 10362
rect 4450 10310 4502 10362
rect 4514 10310 4566 10362
rect 4578 10310 4630 10362
rect 3976 10183 4028 10192
rect 3976 10149 3985 10183
rect 3985 10149 4019 10183
rect 4019 10149 4028 10183
rect 3976 10140 4028 10149
rect 4252 10072 4304 10124
rect 6368 10208 6420 10260
rect 4804 10183 4856 10192
rect 4804 10149 4813 10183
rect 4813 10149 4847 10183
rect 4847 10149 4856 10183
rect 4804 10140 4856 10149
rect 5080 10183 5132 10192
rect 5080 10149 5089 10183
rect 5089 10149 5123 10183
rect 5123 10149 5132 10183
rect 5080 10140 5132 10149
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 5264 10072 5316 10081
rect 5632 10072 5684 10124
rect 5356 10004 5408 10056
rect 5816 10004 5868 10056
rect 4988 9911 5040 9920
rect 4988 9877 4997 9911
rect 4997 9877 5031 9911
rect 5031 9877 5040 9911
rect 4988 9868 5040 9877
rect 5632 9911 5684 9920
rect 5632 9877 5641 9911
rect 5641 9877 5675 9911
rect 5675 9877 5684 9911
rect 5632 9868 5684 9877
rect 9312 10140 9364 10192
rect 16396 10251 16448 10260
rect 16396 10217 16405 10251
rect 16405 10217 16439 10251
rect 16439 10217 16448 10251
rect 16396 10208 16448 10217
rect 6920 10115 6972 10124
rect 6920 10081 6938 10115
rect 6938 10081 6972 10115
rect 6920 10072 6972 10081
rect 8668 10072 8720 10124
rect 8760 10115 8812 10124
rect 8760 10081 8769 10115
rect 8769 10081 8803 10115
rect 8803 10081 8812 10115
rect 8760 10072 8812 10081
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 11704 10115 11756 10124
rect 11704 10081 11713 10115
rect 11713 10081 11747 10115
rect 11747 10081 11756 10115
rect 11704 10072 11756 10081
rect 12440 10115 12492 10124
rect 12440 10081 12449 10115
rect 12449 10081 12483 10115
rect 12483 10081 12492 10115
rect 12440 10072 12492 10081
rect 13820 10115 13872 10124
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 13820 10072 13872 10081
rect 14556 10115 14608 10124
rect 14556 10081 14565 10115
rect 14565 10081 14599 10115
rect 14599 10081 14608 10115
rect 14556 10072 14608 10081
rect 15384 10072 15436 10124
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 17040 10208 17092 10260
rect 17776 10208 17828 10260
rect 21456 10208 21508 10260
rect 22008 10208 22060 10260
rect 22192 10208 22244 10260
rect 21088 10183 21140 10192
rect 21088 10149 21097 10183
rect 21097 10149 21131 10183
rect 21131 10149 21140 10183
rect 21088 10140 21140 10149
rect 17500 10072 17552 10124
rect 18144 10072 18196 10124
rect 20260 10072 20312 10124
rect 8852 10047 8904 10056
rect 8852 10013 8861 10047
rect 8861 10013 8895 10047
rect 8895 10013 8904 10047
rect 8852 10004 8904 10013
rect 11612 10047 11664 10056
rect 11612 10013 11621 10047
rect 11621 10013 11655 10047
rect 11655 10013 11664 10047
rect 11612 10004 11664 10013
rect 12256 10047 12308 10056
rect 12256 10013 12265 10047
rect 12265 10013 12299 10047
rect 12299 10013 12308 10047
rect 12256 10004 12308 10013
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 14740 10004 14792 10056
rect 15108 10047 15160 10056
rect 15108 10013 15117 10047
rect 15117 10013 15151 10047
rect 15151 10013 15160 10047
rect 15108 10004 15160 10013
rect 19892 10047 19944 10056
rect 19892 10013 19901 10047
rect 19901 10013 19935 10047
rect 19935 10013 19944 10047
rect 20812 10115 20864 10124
rect 20812 10081 20821 10115
rect 20821 10081 20855 10115
rect 20855 10081 20864 10115
rect 20812 10072 20864 10081
rect 20904 10115 20956 10124
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 19892 10004 19944 10013
rect 21548 10047 21600 10056
rect 21548 10013 21557 10047
rect 21557 10013 21591 10047
rect 21591 10013 21600 10047
rect 21548 10004 21600 10013
rect 22468 10115 22520 10124
rect 22468 10081 22477 10115
rect 22477 10081 22511 10115
rect 22511 10081 22520 10115
rect 22468 10072 22520 10081
rect 22652 10072 22704 10124
rect 15200 9936 15252 9988
rect 22836 9936 22888 9988
rect 6460 9868 6512 9920
rect 10416 9868 10468 9920
rect 14740 9868 14792 9920
rect 14832 9911 14884 9920
rect 14832 9877 14841 9911
rect 14841 9877 14875 9911
rect 14875 9877 14884 9911
rect 14832 9868 14884 9877
rect 15292 9868 15344 9920
rect 16764 9911 16816 9920
rect 16764 9877 16773 9911
rect 16773 9877 16807 9911
rect 16807 9877 16816 9911
rect 16764 9868 16816 9877
rect 19616 9868 19668 9920
rect 21824 9868 21876 9920
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 4712 9664 4764 9716
rect 5172 9664 5224 9716
rect 5264 9664 5316 9716
rect 6000 9664 6052 9716
rect 6736 9707 6788 9716
rect 6736 9673 6745 9707
rect 6745 9673 6779 9707
rect 6779 9673 6788 9707
rect 6736 9664 6788 9673
rect 6920 9707 6972 9716
rect 6920 9673 6929 9707
rect 6929 9673 6963 9707
rect 6963 9673 6972 9707
rect 6920 9664 6972 9673
rect 9956 9664 10008 9716
rect 12256 9664 12308 9716
rect 14648 9664 14700 9716
rect 14832 9664 14884 9716
rect 16764 9664 16816 9716
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 14464 9596 14516 9648
rect 16580 9596 16632 9648
rect 16672 9596 16724 9648
rect 17776 9707 17828 9716
rect 17776 9673 17785 9707
rect 17785 9673 17819 9707
rect 17819 9673 17828 9707
rect 17776 9664 17828 9673
rect 18236 9664 18288 9716
rect 18420 9664 18472 9716
rect 19248 9707 19300 9716
rect 19248 9673 19257 9707
rect 19257 9673 19291 9707
rect 19291 9673 19300 9707
rect 19248 9664 19300 9673
rect 17500 9639 17552 9648
rect 17500 9605 17509 9639
rect 17509 9605 17543 9639
rect 17543 9605 17552 9639
rect 17500 9596 17552 9605
rect 4896 9571 4948 9580
rect 4896 9537 4905 9571
rect 4905 9537 4939 9571
rect 4939 9537 4948 9571
rect 4896 9528 4948 9537
rect 10324 9528 10376 9580
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 16396 9528 16448 9580
rect 4988 9460 5040 9512
rect 5632 9460 5684 9512
rect 7656 9460 7708 9512
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 9772 9460 9824 9512
rect 12072 9503 12124 9512
rect 12072 9469 12081 9503
rect 12081 9469 12115 9503
rect 12115 9469 12124 9503
rect 12072 9460 12124 9469
rect 14740 9460 14792 9512
rect 15292 9503 15344 9512
rect 15292 9469 15301 9503
rect 15301 9469 15335 9503
rect 15335 9469 15344 9503
rect 15292 9460 15344 9469
rect 15476 9460 15528 9512
rect 16304 9460 16356 9512
rect 16488 9460 16540 9512
rect 17040 9528 17092 9580
rect 20812 9664 20864 9716
rect 20996 9596 21048 9648
rect 5264 9392 5316 9444
rect 6920 9392 6972 9444
rect 4804 9324 4856 9376
rect 5172 9324 5224 9376
rect 7564 9367 7616 9376
rect 7564 9333 7573 9367
rect 7573 9333 7607 9367
rect 7607 9333 7616 9367
rect 7564 9324 7616 9333
rect 8576 9392 8628 9444
rect 10876 9392 10928 9444
rect 13820 9392 13872 9444
rect 14280 9392 14332 9444
rect 14924 9392 14976 9444
rect 17868 9392 17920 9444
rect 19616 9503 19668 9512
rect 19616 9469 19625 9503
rect 19625 9469 19659 9503
rect 19659 9469 19668 9503
rect 19616 9460 19668 9469
rect 21180 9460 21232 9512
rect 21824 9503 21876 9512
rect 21824 9469 21858 9503
rect 21858 9469 21876 9503
rect 21824 9460 21876 9469
rect 20168 9392 20220 9444
rect 8208 9324 8260 9376
rect 8944 9367 8996 9376
rect 8944 9333 8953 9367
rect 8953 9333 8987 9367
rect 8987 9333 8996 9367
rect 8944 9324 8996 9333
rect 9496 9324 9548 9376
rect 12992 9324 13044 9376
rect 16764 9324 16816 9376
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 18788 9367 18840 9376
rect 18788 9333 18797 9367
rect 18797 9333 18831 9367
rect 18831 9333 18840 9367
rect 18788 9324 18840 9333
rect 19156 9324 19208 9376
rect 19708 9324 19760 9376
rect 19800 9324 19852 9376
rect 19984 9324 20036 9376
rect 20536 9324 20588 9376
rect 22652 9324 22704 9376
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 5264 9163 5316 9172
rect 5264 9129 5273 9163
rect 5273 9129 5307 9163
rect 5307 9129 5316 9163
rect 5264 9120 5316 9129
rect 7564 9120 7616 9172
rect 9772 9120 9824 9172
rect 9956 9163 10008 9172
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 5080 9052 5132 9104
rect 6920 9095 6972 9104
rect 5356 8984 5408 9036
rect 5264 8916 5316 8968
rect 6920 9061 6929 9095
rect 6929 9061 6963 9095
rect 6963 9061 6972 9095
rect 6920 9052 6972 9061
rect 7748 9052 7800 9104
rect 7840 9052 7892 9104
rect 8760 9052 8812 9104
rect 9588 9027 9640 9036
rect 9588 8993 9597 9027
rect 9597 8993 9631 9027
rect 9631 8993 9640 9027
rect 9588 8984 9640 8993
rect 10784 9120 10836 9172
rect 12072 9120 12124 9172
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 10876 8984 10928 9036
rect 11612 9027 11664 9036
rect 11612 8993 11621 9027
rect 11621 8993 11655 9027
rect 11655 8993 11664 9027
rect 11612 8984 11664 8993
rect 13084 9095 13136 9104
rect 13084 9061 13093 9095
rect 13093 9061 13127 9095
rect 13127 9061 13136 9095
rect 13084 9052 13136 9061
rect 12808 8984 12860 9036
rect 7104 8823 7156 8832
rect 7104 8789 7113 8823
rect 7113 8789 7147 8823
rect 7147 8789 7156 8823
rect 7104 8780 7156 8789
rect 8576 8848 8628 8900
rect 9588 8848 9640 8900
rect 10692 8848 10744 8900
rect 8668 8780 8720 8832
rect 10232 8823 10284 8832
rect 10232 8789 10241 8823
rect 10241 8789 10275 8823
rect 10275 8789 10284 8823
rect 10232 8780 10284 8789
rect 10600 8780 10652 8832
rect 11612 8848 11664 8900
rect 13728 8984 13780 9036
rect 14280 8984 14332 9036
rect 15384 9095 15436 9104
rect 15384 9061 15393 9095
rect 15393 9061 15427 9095
rect 15427 9061 15436 9095
rect 15384 9052 15436 9061
rect 14464 9027 14516 9036
rect 14464 8993 14473 9027
rect 14473 8993 14507 9027
rect 14507 8993 14516 9027
rect 14464 8984 14516 8993
rect 14740 9027 14792 9036
rect 14740 8993 14749 9027
rect 14749 8993 14783 9027
rect 14783 8993 14792 9027
rect 14740 8984 14792 8993
rect 14924 9027 14976 9036
rect 14924 8993 14933 9027
rect 14933 8993 14967 9027
rect 14967 8993 14976 9027
rect 14924 8984 14976 8993
rect 15016 8984 15068 9036
rect 11244 8780 11296 8832
rect 12440 8823 12492 8832
rect 12440 8789 12449 8823
rect 12449 8789 12483 8823
rect 12483 8789 12492 8823
rect 12440 8780 12492 8789
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 13912 8823 13964 8832
rect 13912 8789 13921 8823
rect 13921 8789 13955 8823
rect 13955 8789 13964 8823
rect 13912 8780 13964 8789
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 15384 8916 15436 8968
rect 15108 8891 15160 8900
rect 15108 8857 15117 8891
rect 15117 8857 15151 8891
rect 15151 8857 15160 8891
rect 15108 8848 15160 8857
rect 15476 8848 15528 8900
rect 15200 8780 15252 8832
rect 15292 8780 15344 8832
rect 17592 9027 17644 9036
rect 18144 9052 18196 9104
rect 18236 9095 18288 9104
rect 18236 9061 18245 9095
rect 18245 9061 18279 9095
rect 18279 9061 18288 9095
rect 18236 9052 18288 9061
rect 18788 9120 18840 9172
rect 20168 9163 20220 9172
rect 20168 9129 20177 9163
rect 20177 9129 20211 9163
rect 20211 9129 20220 9163
rect 20168 9120 20220 9129
rect 22560 9120 22612 9172
rect 20076 9052 20128 9104
rect 20444 9052 20496 9104
rect 20536 9052 20588 9104
rect 17592 8993 17610 9027
rect 17610 8993 17644 9027
rect 17592 8984 17644 8993
rect 16396 8848 16448 8900
rect 19248 8984 19300 9036
rect 20168 8984 20220 9036
rect 20260 8984 20312 9036
rect 20628 8984 20680 9036
rect 21272 9052 21324 9104
rect 22744 8984 22796 9036
rect 18328 8780 18380 8832
rect 18420 8823 18472 8832
rect 18420 8789 18429 8823
rect 18429 8789 18463 8823
rect 18463 8789 18472 8823
rect 18420 8780 18472 8789
rect 18880 8780 18932 8832
rect 21180 8916 21232 8968
rect 21364 8959 21416 8968
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 19800 8848 19852 8900
rect 20168 8780 20220 8832
rect 20720 8780 20772 8832
rect 20996 8780 21048 8832
rect 21548 8780 21600 8832
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 7104 8576 7156 8628
rect 7840 8576 7892 8628
rect 8392 8576 8444 8628
rect 9772 8576 9824 8628
rect 10324 8619 10376 8628
rect 10324 8585 10333 8619
rect 10333 8585 10367 8619
rect 10367 8585 10376 8619
rect 10324 8576 10376 8585
rect 12440 8576 12492 8628
rect 12808 8619 12860 8628
rect 12808 8585 12817 8619
rect 12817 8585 12851 8619
rect 12851 8585 12860 8619
rect 12808 8576 12860 8585
rect 4896 8508 4948 8560
rect 8300 8508 8352 8560
rect 11060 8508 11112 8560
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 11244 8440 11296 8492
rect 5632 8372 5684 8424
rect 7656 8372 7708 8424
rect 4712 8236 4764 8288
rect 7472 8304 7524 8356
rect 6000 8236 6052 8288
rect 6920 8236 6972 8288
rect 8484 8372 8536 8424
rect 8668 8372 8720 8424
rect 11336 8372 11388 8424
rect 9312 8304 9364 8356
rect 10140 8304 10192 8356
rect 12992 8347 13044 8356
rect 12992 8313 13001 8347
rect 13001 8313 13035 8347
rect 13035 8313 13044 8347
rect 12992 8304 13044 8313
rect 13452 8304 13504 8356
rect 13728 8415 13780 8424
rect 13728 8381 13737 8415
rect 13737 8381 13771 8415
rect 13771 8381 13780 8415
rect 13728 8372 13780 8381
rect 15016 8576 15068 8628
rect 15384 8576 15436 8628
rect 16396 8576 16448 8628
rect 13912 8372 13964 8424
rect 15016 8372 15068 8424
rect 16856 8576 16908 8628
rect 17592 8619 17644 8628
rect 17592 8585 17601 8619
rect 17601 8585 17635 8619
rect 17635 8585 17644 8619
rect 17592 8576 17644 8585
rect 18328 8576 18380 8628
rect 19984 8576 20036 8628
rect 20444 8619 20496 8628
rect 20444 8585 20453 8619
rect 20453 8585 20487 8619
rect 20487 8585 20496 8619
rect 20444 8576 20496 8585
rect 22376 8576 22428 8628
rect 22560 8576 22612 8628
rect 19892 8508 19944 8560
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 19156 8415 19208 8424
rect 14924 8304 14976 8356
rect 15476 8304 15528 8356
rect 16580 8304 16632 8356
rect 17224 8347 17276 8356
rect 13360 8279 13412 8288
rect 13360 8245 13369 8279
rect 13369 8245 13403 8279
rect 13403 8245 13412 8279
rect 13360 8236 13412 8245
rect 14280 8236 14332 8288
rect 14740 8236 14792 8288
rect 15384 8236 15436 8288
rect 17224 8313 17233 8347
rect 17233 8313 17267 8347
rect 17267 8313 17276 8347
rect 17224 8304 17276 8313
rect 19156 8381 19190 8415
rect 19190 8381 19208 8415
rect 19156 8372 19208 8381
rect 20812 8508 20864 8560
rect 20720 8304 20772 8356
rect 20996 8415 21048 8424
rect 20996 8381 21005 8415
rect 21005 8381 21039 8415
rect 21039 8381 21048 8415
rect 20996 8372 21048 8381
rect 21180 8415 21232 8424
rect 21180 8381 21189 8415
rect 21189 8381 21223 8415
rect 21223 8381 21232 8415
rect 21180 8372 21232 8381
rect 21916 8508 21968 8560
rect 22744 8551 22796 8560
rect 22744 8517 22753 8551
rect 22753 8517 22787 8551
rect 22787 8517 22796 8551
rect 22744 8508 22796 8517
rect 21456 8440 21508 8492
rect 21640 8483 21692 8492
rect 21640 8449 21649 8483
rect 21649 8449 21683 8483
rect 21683 8449 21692 8483
rect 21640 8440 21692 8449
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 22008 8415 22060 8424
rect 22008 8381 22017 8415
rect 22017 8381 22051 8415
rect 22051 8381 22060 8415
rect 22008 8372 22060 8381
rect 22928 8415 22980 8424
rect 22928 8381 22937 8415
rect 22937 8381 22971 8415
rect 22971 8381 22980 8415
rect 22928 8372 22980 8381
rect 21548 8304 21600 8356
rect 22192 8304 22244 8356
rect 22652 8347 22704 8356
rect 22652 8313 22661 8347
rect 22661 8313 22695 8347
rect 22695 8313 22704 8347
rect 22652 8304 22704 8313
rect 20904 8236 20956 8288
rect 21456 8236 21508 8288
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 5908 8032 5960 8084
rect 7840 8075 7892 8084
rect 7840 8041 7849 8075
rect 7849 8041 7883 8075
rect 7883 8041 7892 8075
rect 7840 8032 7892 8041
rect 8208 8032 8260 8084
rect 4436 7964 4488 8016
rect 8944 8007 8996 8016
rect 8944 7973 8962 8007
rect 8962 7973 8996 8007
rect 9312 8075 9364 8084
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 10324 8075 10376 8084
rect 10324 8041 10333 8075
rect 10333 8041 10367 8075
rect 10367 8041 10376 8075
rect 10324 8032 10376 8041
rect 8944 7964 8996 7973
rect 10140 8007 10192 8016
rect 10140 7973 10149 8007
rect 10149 7973 10183 8007
rect 10183 7973 10192 8007
rect 10140 7964 10192 7973
rect 4528 7896 4580 7948
rect 5080 7828 5132 7880
rect 4988 7760 5040 7812
rect 5264 7803 5316 7812
rect 5264 7769 5273 7803
rect 5273 7769 5307 7803
rect 5307 7769 5316 7803
rect 5264 7760 5316 7769
rect 5172 7735 5224 7744
rect 5172 7701 5181 7735
rect 5181 7701 5215 7735
rect 5215 7701 5224 7735
rect 5172 7692 5224 7701
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 6276 7828 6328 7837
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 7104 7896 7156 7948
rect 8668 7896 8720 7948
rect 11612 8032 11664 8084
rect 13820 8032 13872 8084
rect 14464 8032 14516 8084
rect 15200 8032 15252 8084
rect 15384 8032 15436 8084
rect 15476 8075 15528 8084
rect 15476 8041 15485 8075
rect 15485 8041 15519 8075
rect 15519 8041 15528 8075
rect 15476 8032 15528 8041
rect 18420 8032 18472 8084
rect 19708 8075 19760 8084
rect 19708 8041 19717 8075
rect 19717 8041 19751 8075
rect 19751 8041 19760 8075
rect 19708 8032 19760 8041
rect 20628 8075 20680 8084
rect 10876 7964 10928 8016
rect 11060 7964 11112 8016
rect 11336 7964 11388 8016
rect 10784 7939 10836 7948
rect 10784 7905 10793 7939
rect 10793 7905 10827 7939
rect 10827 7905 10836 7939
rect 10784 7896 10836 7905
rect 13084 7939 13136 7948
rect 13084 7905 13093 7939
rect 13093 7905 13127 7939
rect 13127 7905 13136 7939
rect 13084 7896 13136 7905
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 13360 7964 13412 8016
rect 19616 8007 19668 8016
rect 19616 7973 19625 8007
rect 19625 7973 19659 8007
rect 19659 7973 19668 8007
rect 19616 7964 19668 7973
rect 19892 8007 19944 8016
rect 19892 7973 19901 8007
rect 19901 7973 19935 8007
rect 19935 7973 19944 8007
rect 19892 7964 19944 7973
rect 20628 8041 20637 8075
rect 20637 8041 20671 8075
rect 20671 8041 20680 8075
rect 20628 8032 20680 8041
rect 20720 7964 20772 8016
rect 21916 8032 21968 8084
rect 22008 8032 22060 8084
rect 15108 7896 15160 7948
rect 19800 7896 19852 7948
rect 20904 7964 20956 8016
rect 21640 7964 21692 8016
rect 21364 7896 21416 7948
rect 6920 7760 6972 7812
rect 6828 7692 6880 7744
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 15292 7735 15344 7744
rect 15292 7701 15301 7735
rect 15301 7701 15335 7735
rect 15335 7701 15344 7735
rect 15292 7692 15344 7701
rect 20812 7735 20864 7744
rect 20812 7701 20821 7735
rect 20821 7701 20855 7735
rect 20855 7701 20864 7735
rect 20812 7692 20864 7701
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 4436 7531 4488 7540
rect 4436 7497 4445 7531
rect 4445 7497 4479 7531
rect 4479 7497 4488 7531
rect 4436 7488 4488 7497
rect 4988 7531 5040 7540
rect 4988 7497 4997 7531
rect 4997 7497 5031 7531
rect 5031 7497 5040 7531
rect 4988 7488 5040 7497
rect 6276 7488 6328 7540
rect 4252 7327 4304 7336
rect 4252 7293 4261 7327
rect 4261 7293 4295 7327
rect 4295 7293 4304 7327
rect 4252 7284 4304 7293
rect 4528 7327 4580 7336
rect 4528 7293 4537 7327
rect 4537 7293 4571 7327
rect 4571 7293 4580 7327
rect 4528 7284 4580 7293
rect 5264 7327 5316 7336
rect 5264 7293 5273 7327
rect 5273 7293 5307 7327
rect 5307 7293 5316 7327
rect 5264 7284 5316 7293
rect 5356 7284 5408 7336
rect 8208 7488 8260 7540
rect 10876 7488 10928 7540
rect 14096 7531 14148 7540
rect 14096 7497 14105 7531
rect 14105 7497 14139 7531
rect 14139 7497 14148 7531
rect 14096 7488 14148 7497
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 6828 7420 6880 7472
rect 8668 7463 8720 7472
rect 8668 7429 8677 7463
rect 8677 7429 8711 7463
rect 8711 7429 8720 7463
rect 8668 7420 8720 7429
rect 4712 7216 4764 7268
rect 5080 7216 5132 7268
rect 7104 7327 7156 7336
rect 7104 7293 7113 7327
rect 7113 7293 7147 7327
rect 7147 7293 7156 7327
rect 7104 7284 7156 7293
rect 8300 7284 8352 7336
rect 11060 7284 11112 7336
rect 14280 7327 14332 7336
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 14464 7327 14516 7336
rect 14464 7293 14473 7327
rect 14473 7293 14507 7327
rect 14507 7293 14516 7327
rect 14464 7284 14516 7293
rect 14924 7284 14976 7336
rect 20904 7284 20956 7336
rect 21916 7284 21968 7336
rect 6920 7259 6972 7268
rect 6920 7225 6929 7259
rect 6929 7225 6963 7259
rect 6963 7225 6972 7259
rect 6920 7216 6972 7225
rect 7472 7216 7524 7268
rect 7748 7259 7800 7268
rect 7748 7225 7757 7259
rect 7757 7225 7791 7259
rect 7791 7225 7800 7259
rect 7748 7216 7800 7225
rect 7380 7191 7432 7200
rect 7380 7157 7389 7191
rect 7389 7157 7423 7191
rect 7423 7157 7432 7191
rect 7380 7148 7432 7157
rect 10416 7148 10468 7200
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 4252 6987 4304 6996
rect 4252 6953 4261 6987
rect 4261 6953 4295 6987
rect 4295 6953 4304 6987
rect 4252 6944 4304 6953
rect 5632 6944 5684 6996
rect 6920 6944 6972 6996
rect 7748 6944 7800 6996
rect 10416 6987 10468 6996
rect 10416 6953 10425 6987
rect 10425 6953 10459 6987
rect 10459 6953 10468 6987
rect 10416 6944 10468 6953
rect 10600 6987 10652 6996
rect 10600 6953 10627 6987
rect 10627 6953 10652 6987
rect 10600 6944 10652 6953
rect 5172 6876 5224 6928
rect 6828 6876 6880 6928
rect 5908 6808 5960 6860
rect 7104 6808 7156 6860
rect 10140 6876 10192 6928
rect 5816 6783 5868 6792
rect 5264 6604 5316 6656
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 10232 6604 10284 6656
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 4712 6400 4764 6452
rect 5816 6400 5868 6452
rect 8668 6264 8720 6316
rect 7380 6128 7432 6180
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 22928 4224 22980 4276
rect 23020 4063 23072 4072
rect 23020 4029 23029 4063
rect 23029 4029 23063 4063
rect 23063 4029 23072 4063
rect 23020 4020 23072 4029
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
<< metal2 >>
rect 1674 23746 1730 24000
rect 4618 23746 4674 24000
rect 1674 23718 1808 23746
rect 1674 23600 1730 23718
rect 1780 23186 1808 23718
rect 4618 23718 4752 23746
rect 4618 23600 4674 23718
rect 4322 23420 4630 23429
rect 4322 23418 4328 23420
rect 4384 23418 4408 23420
rect 4464 23418 4488 23420
rect 4544 23418 4568 23420
rect 4624 23418 4630 23420
rect 4384 23366 4386 23418
rect 4566 23366 4568 23418
rect 4322 23364 4328 23366
rect 4384 23364 4408 23366
rect 4464 23364 4488 23366
rect 4544 23364 4568 23366
rect 4624 23364 4630 23366
rect 4322 23355 4630 23364
rect 4724 23186 4752 23718
rect 7562 23600 7618 24000
rect 10506 23746 10562 24000
rect 10428 23718 10562 23746
rect 7576 23322 7604 23600
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7656 23316 7708 23322
rect 7656 23258 7708 23264
rect 1768 23180 1820 23186
rect 1768 23122 1820 23128
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 6276 23180 6328 23186
rect 6276 23122 6328 23128
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 5448 23044 5500 23050
rect 5448 22986 5500 22992
rect 6184 23044 6236 23050
rect 6184 22986 6236 22992
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 5356 22976 5408 22982
rect 5356 22918 5408 22924
rect 3662 22876 3970 22885
rect 3662 22874 3668 22876
rect 3724 22874 3748 22876
rect 3804 22874 3828 22876
rect 3884 22874 3908 22876
rect 3964 22874 3970 22876
rect 3724 22822 3726 22874
rect 3906 22822 3908 22874
rect 3662 22820 3668 22822
rect 3724 22820 3748 22822
rect 3804 22820 3828 22822
rect 3884 22820 3908 22822
rect 3964 22820 3970 22822
rect 3662 22811 3970 22820
rect 4908 22642 4936 22918
rect 5368 22710 5396 22918
rect 5356 22704 5408 22710
rect 5356 22646 5408 22652
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 4908 22506 4936 22578
rect 4896 22500 4948 22506
rect 4896 22442 4948 22448
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 4322 22332 4630 22341
rect 4322 22330 4328 22332
rect 4384 22330 4408 22332
rect 4464 22330 4488 22332
rect 4544 22330 4568 22332
rect 4624 22330 4630 22332
rect 4384 22278 4386 22330
rect 4566 22278 4568 22330
rect 4322 22276 4328 22278
rect 4384 22276 4408 22278
rect 4464 22276 4488 22278
rect 4544 22276 4568 22278
rect 4624 22276 4630 22278
rect 4322 22267 4630 22276
rect 3662 21788 3970 21797
rect 3662 21786 3668 21788
rect 3724 21786 3748 21788
rect 3804 21786 3828 21788
rect 3884 21786 3908 21788
rect 3964 21786 3970 21788
rect 3724 21734 3726 21786
rect 3906 21734 3908 21786
rect 3662 21732 3668 21734
rect 3724 21732 3748 21734
rect 3804 21732 3828 21734
rect 3884 21732 3908 21734
rect 3964 21732 3970 21734
rect 3662 21723 3970 21732
rect 4712 21616 4764 21622
rect 4712 21558 4764 21564
rect 4322 21244 4630 21253
rect 4322 21242 4328 21244
rect 4384 21242 4408 21244
rect 4464 21242 4488 21244
rect 4544 21242 4568 21244
rect 4624 21242 4630 21244
rect 4384 21190 4386 21242
rect 4566 21190 4568 21242
rect 4322 21188 4328 21190
rect 4384 21188 4408 21190
rect 4464 21188 4488 21190
rect 4544 21188 4568 21190
rect 4624 21188 4630 21190
rect 4322 21179 4630 21188
rect 4724 21026 4752 21558
rect 5092 21418 5120 22374
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 5276 21622 5304 21830
rect 5264 21616 5316 21622
rect 5264 21558 5316 21564
rect 5080 21412 5132 21418
rect 5080 21354 5132 21360
rect 5264 21412 5316 21418
rect 5264 21354 5316 21360
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 5184 21078 5212 21286
rect 4632 20998 4752 21026
rect 5172 21072 5224 21078
rect 5172 21014 5224 21020
rect 4632 20942 4660 20998
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 3662 20700 3970 20709
rect 3662 20698 3668 20700
rect 3724 20698 3748 20700
rect 3804 20698 3828 20700
rect 3884 20698 3908 20700
rect 3964 20698 3970 20700
rect 3724 20646 3726 20698
rect 3906 20646 3908 20698
rect 3662 20644 3668 20646
rect 3724 20644 3748 20646
rect 3804 20644 3828 20646
rect 3884 20644 3908 20646
rect 3964 20644 3970 20646
rect 3662 20635 3970 20644
rect 4322 20156 4630 20165
rect 4322 20154 4328 20156
rect 4384 20154 4408 20156
rect 4464 20154 4488 20156
rect 4544 20154 4568 20156
rect 4624 20154 4630 20156
rect 4384 20102 4386 20154
rect 4566 20102 4568 20154
rect 4322 20100 4328 20102
rect 4384 20100 4408 20102
rect 4464 20100 4488 20102
rect 4544 20100 4568 20102
rect 4624 20100 4630 20102
rect 4322 20091 4630 20100
rect 3662 19612 3970 19621
rect 3662 19610 3668 19612
rect 3724 19610 3748 19612
rect 3804 19610 3828 19612
rect 3884 19610 3908 19612
rect 3964 19610 3970 19612
rect 3724 19558 3726 19610
rect 3906 19558 3908 19610
rect 3662 19556 3668 19558
rect 3724 19556 3748 19558
rect 3804 19556 3828 19558
rect 3884 19556 3908 19558
rect 3964 19556 3970 19558
rect 3662 19547 3970 19556
rect 4724 19242 4752 20998
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 5092 20806 5120 20878
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 5092 20602 5120 20742
rect 5080 20596 5132 20602
rect 5080 20538 5132 20544
rect 5184 20466 5212 21014
rect 5276 21010 5304 21354
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5172 20460 5224 20466
rect 5172 20402 5224 20408
rect 4712 19236 4764 19242
rect 4712 19178 4764 19184
rect 5276 19174 5304 20946
rect 5368 20874 5396 22646
rect 5460 22574 5488 22986
rect 5632 22636 5684 22642
rect 5632 22578 5684 22584
rect 5448 22568 5500 22574
rect 5448 22510 5500 22516
rect 5460 22438 5488 22510
rect 5448 22432 5500 22438
rect 5448 22374 5500 22380
rect 5644 22098 5672 22578
rect 6196 22506 6224 22986
rect 6000 22500 6052 22506
rect 6000 22442 6052 22448
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 5632 22092 5684 22098
rect 5632 22034 5684 22040
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 5644 21010 5672 21082
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5356 20868 5408 20874
rect 5356 20810 5408 20816
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 4322 19068 4630 19077
rect 4322 19066 4328 19068
rect 4384 19066 4408 19068
rect 4464 19066 4488 19068
rect 4544 19066 4568 19068
rect 4624 19066 4630 19068
rect 4384 19014 4386 19066
rect 4566 19014 4568 19066
rect 4322 19012 4328 19014
rect 4384 19012 4408 19014
rect 4464 19012 4488 19014
rect 4544 19012 4568 19014
rect 4624 19012 4630 19014
rect 4322 19003 4630 19012
rect 5276 18698 5304 19110
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 3662 18459 3970 18468
rect 5276 18290 5304 18634
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 4804 18216 4856 18222
rect 5276 18170 5304 18226
rect 4804 18158 4856 18164
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4322 17980 4630 17989
rect 4322 17978 4328 17980
rect 4384 17978 4408 17980
rect 4464 17978 4488 17980
rect 4544 17978 4568 17980
rect 4624 17978 4630 17980
rect 4384 17926 4386 17978
rect 4566 17926 4568 17978
rect 4322 17924 4328 17926
rect 4384 17924 4408 17926
rect 4464 17924 4488 17926
rect 4544 17924 4568 17926
rect 4624 17924 4630 17926
rect 4322 17915 4630 17924
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 4322 16892 4630 16901
rect 4322 16890 4328 16892
rect 4384 16890 4408 16892
rect 4464 16890 4488 16892
rect 4544 16890 4568 16892
rect 4624 16890 4630 16892
rect 4384 16838 4386 16890
rect 4566 16838 4568 16890
rect 4322 16836 4328 16838
rect 4384 16836 4408 16838
rect 4464 16836 4488 16838
rect 4544 16836 4568 16838
rect 4624 16836 4630 16838
rect 4322 16827 4630 16836
rect 4724 16658 4752 18090
rect 4816 17814 4844 18158
rect 5184 18142 5304 18170
rect 5368 18154 5396 20810
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5460 20602 5488 20742
rect 5448 20596 5500 20602
rect 5448 20538 5500 20544
rect 5460 20398 5488 20538
rect 5644 20466 5672 20946
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5908 20460 5960 20466
rect 5908 20402 5960 20408
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 5460 18834 5488 19178
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5460 18222 5488 18770
rect 5552 18766 5580 19858
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5356 18148 5408 18154
rect 5184 17882 5212 18142
rect 5356 18090 5408 18096
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 4804 17808 4856 17814
rect 4804 17750 4856 17756
rect 4816 16658 4844 17750
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4908 16794 4936 17070
rect 5184 16998 5212 17818
rect 5264 17808 5316 17814
rect 5460 17762 5488 18158
rect 5552 17882 5580 18702
rect 5644 18426 5672 19450
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5264 17750 5316 17756
rect 5276 17134 5304 17750
rect 5368 17746 5488 17762
rect 5644 17746 5672 18362
rect 5356 17740 5488 17746
rect 5408 17734 5488 17740
rect 5356 17682 5408 17688
rect 5460 17542 5488 17734
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5552 17218 5580 17614
rect 5368 17190 5580 17218
rect 5368 17134 5396 17190
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 4816 15978 4844 16594
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4322 15804 4630 15813
rect 4322 15802 4328 15804
rect 4384 15802 4408 15804
rect 4464 15802 4488 15804
rect 4544 15802 4568 15804
rect 4624 15802 4630 15804
rect 4384 15750 4386 15802
rect 4566 15750 4568 15802
rect 4322 15748 4328 15750
rect 4384 15748 4408 15750
rect 4464 15748 4488 15750
rect 4544 15748 4568 15750
rect 4624 15748 4630 15750
rect 4322 15739 4630 15748
rect 4908 15638 4936 16730
rect 5460 16726 5488 17070
rect 5448 16720 5500 16726
rect 5448 16662 5500 16668
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5080 16176 5132 16182
rect 5080 16118 5132 16124
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 5092 15570 5120 16118
rect 5552 16046 5580 16526
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5644 15570 5672 15914
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 4322 14716 4630 14725
rect 4322 14714 4328 14716
rect 4384 14714 4408 14716
rect 4464 14714 4488 14716
rect 4544 14714 4568 14716
rect 4624 14714 4630 14716
rect 4384 14662 4386 14714
rect 4566 14662 4568 14714
rect 4322 14660 4328 14662
rect 4384 14660 4408 14662
rect 4464 14660 4488 14662
rect 4544 14660 4568 14662
rect 4624 14660 4630 14662
rect 4322 14651 4630 14660
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 4322 13628 4630 13637
rect 4322 13626 4328 13628
rect 4384 13626 4408 13628
rect 4464 13626 4488 13628
rect 4544 13626 4568 13628
rect 4624 13626 4630 13628
rect 4384 13574 4386 13626
rect 4566 13574 4568 13626
rect 4322 13572 4328 13574
rect 4384 13572 4408 13574
rect 4464 13572 4488 13574
rect 4544 13572 4568 13574
rect 4624 13572 4630 13574
rect 4322 13563 4630 13572
rect 5552 13530 5580 13806
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5736 13462 5764 20198
rect 5920 17270 5948 20402
rect 6012 20398 6040 22442
rect 6196 21554 6224 22442
rect 6288 22098 6316 23122
rect 6920 23112 6972 23118
rect 6920 23054 6972 23060
rect 6368 22568 6420 22574
rect 6368 22510 6420 22516
rect 6276 22092 6328 22098
rect 6276 22034 6328 22040
rect 6380 21894 6408 22510
rect 6932 22098 6960 23054
rect 7392 22710 7420 23122
rect 7668 23118 7696 23258
rect 10428 23254 10456 23718
rect 10506 23600 10562 23718
rect 13450 23746 13506 24000
rect 13450 23718 13584 23746
rect 13450 23600 13506 23718
rect 10416 23248 10468 23254
rect 10416 23190 10468 23196
rect 13556 23186 13584 23718
rect 16394 23600 16450 24000
rect 19338 23746 19394 24000
rect 19338 23718 19564 23746
rect 19338 23600 19394 23718
rect 14464 23248 14516 23254
rect 14464 23190 14516 23196
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 7656 23112 7708 23118
rect 7656 23054 7708 23060
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7380 22704 7432 22710
rect 7380 22646 7432 22652
rect 7196 22568 7248 22574
rect 7196 22510 7248 22516
rect 6920 22092 6972 22098
rect 6920 22034 6972 22040
rect 6368 21888 6420 21894
rect 6368 21830 6420 21836
rect 6380 21554 6408 21830
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 6368 21548 6420 21554
rect 6368 21490 6420 21496
rect 6368 21412 6420 21418
rect 6368 21354 6420 21360
rect 6380 21146 6408 21354
rect 6368 21140 6420 21146
rect 6368 21082 6420 21088
rect 6932 21010 6960 22034
rect 7208 21554 7236 22510
rect 7392 21962 7420 22646
rect 7656 22500 7708 22506
rect 7656 22442 7708 22448
rect 7564 22160 7616 22166
rect 7564 22102 7616 22108
rect 7380 21956 7432 21962
rect 7380 21898 7432 21904
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7484 21554 7512 21898
rect 7576 21706 7604 22102
rect 7668 21962 7696 22442
rect 7656 21956 7708 21962
rect 7656 21898 7708 21904
rect 7576 21678 7696 21706
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 7472 21548 7524 21554
rect 7472 21490 7524 21496
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 6000 20392 6052 20398
rect 6104 20380 6132 20538
rect 6656 20398 6684 20742
rect 7116 20398 7144 20946
rect 6052 20352 6132 20380
rect 6000 20334 6052 20340
rect 6000 19984 6052 19990
rect 6000 19926 6052 19932
rect 6012 18970 6040 19926
rect 6104 19922 6132 20352
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7380 20324 7432 20330
rect 7380 20266 7432 20272
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 6012 18222 6040 18906
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 6012 17678 6040 18158
rect 6288 18086 6316 18770
rect 6380 18154 6408 20198
rect 6932 19922 6960 20198
rect 7392 20058 7420 20266
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6840 19310 6868 19722
rect 6932 19310 6960 19858
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 6644 18760 6696 18766
rect 6642 18728 6644 18737
rect 6696 18728 6698 18737
rect 6642 18663 6698 18672
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6748 18290 6776 18566
rect 6840 18426 6868 18770
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 7208 18290 7236 18770
rect 7300 18290 7328 19110
rect 7484 18834 7512 21490
rect 7576 20074 7604 21558
rect 7668 21418 7696 21678
rect 7760 21486 7788 22918
rect 9232 22574 9260 23122
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 10968 23112 11020 23118
rect 10968 23054 11020 23060
rect 9404 23044 9456 23050
rect 9404 22986 9456 22992
rect 9416 22642 9444 22986
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9220 22568 9272 22574
rect 9220 22510 9272 22516
rect 8484 22432 8536 22438
rect 8484 22374 8536 22380
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 8220 21962 8248 22034
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 7748 21480 7800 21486
rect 7748 21422 7800 21428
rect 8220 21418 8248 21898
rect 8496 21554 8524 22374
rect 9048 21690 9076 22374
rect 9232 22166 9260 22510
rect 9220 22160 9272 22166
rect 9220 22102 9272 22108
rect 9220 22024 9272 22030
rect 9220 21966 9272 21972
rect 9036 21684 9088 21690
rect 9036 21626 9088 21632
rect 9232 21554 9260 21966
rect 9416 21894 9444 22578
rect 9600 22506 9628 23054
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 10416 22772 10468 22778
rect 10416 22714 10468 22720
rect 9784 22506 9812 22714
rect 9956 22704 10008 22710
rect 9956 22646 10008 22652
rect 9588 22500 9640 22506
rect 9588 22442 9640 22448
rect 9772 22500 9824 22506
rect 9772 22442 9824 22448
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 7656 21412 7708 21418
rect 7656 21354 7708 21360
rect 8116 21412 8168 21418
rect 8116 21354 8168 21360
rect 8208 21412 8260 21418
rect 8208 21354 8260 21360
rect 8128 21146 8156 21354
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 7932 21072 7984 21078
rect 7932 21014 7984 21020
rect 7944 20398 7972 21014
rect 8220 21010 8248 21354
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7576 20046 7696 20074
rect 7944 20058 7972 20334
rect 7564 19916 7616 19922
rect 7564 19858 7616 19864
rect 7576 19514 7604 19858
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7576 18970 7604 19178
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7024 18170 7052 18226
rect 6368 18148 6420 18154
rect 7024 18142 7144 18170
rect 6368 18090 6420 18096
rect 7116 18086 7144 18142
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 6288 17746 6316 18022
rect 6564 17746 6592 18022
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 6012 17338 6040 17614
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 6368 17264 6420 17270
rect 6368 17206 6420 17212
rect 5816 17060 5868 17066
rect 5816 17002 5868 17008
rect 5828 16590 5856 17002
rect 5920 16658 5948 17206
rect 6380 17134 6408 17206
rect 6472 17134 6500 17478
rect 6564 17134 6592 17682
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6368 17128 6420 17134
rect 6368 17070 6420 17076
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 6104 16590 6132 16934
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6460 16516 6512 16522
rect 6460 16458 6512 16464
rect 6472 16046 6500 16458
rect 6932 16114 6960 17274
rect 7024 17134 7052 17614
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 7116 16658 7144 18022
rect 7208 17678 7236 18226
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7484 16726 7512 18770
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7116 16250 7144 16594
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7208 16114 7236 16390
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5828 13734 5856 15438
rect 6196 14618 6224 15982
rect 7484 15570 7512 16118
rect 7576 16046 7604 18906
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7576 15706 7604 15982
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 7472 15564 7524 15570
rect 7472 15506 7524 15512
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6380 14414 6408 15506
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5724 13456 5776 13462
rect 5724 13398 5776 13404
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 6012 12782 6040 14214
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6196 13530 6224 14010
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 6196 12714 6224 13466
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6184 12708 6236 12714
rect 6184 12650 6236 12656
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 4322 12540 4630 12549
rect 4322 12538 4328 12540
rect 4384 12538 4408 12540
rect 4464 12538 4488 12540
rect 4544 12538 4568 12540
rect 4624 12538 4630 12540
rect 4384 12486 4386 12538
rect 4566 12486 4568 12538
rect 4322 12484 4328 12486
rect 4384 12484 4408 12486
rect 4464 12484 4488 12486
rect 4544 12484 4568 12486
rect 4624 12484 4630 12486
rect 4322 12475 4630 12484
rect 5552 12374 5580 12582
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 4322 11452 4630 11461
rect 4322 11450 4328 11452
rect 4384 11450 4408 11452
rect 4464 11450 4488 11452
rect 4544 11450 4568 11452
rect 4624 11450 4630 11452
rect 4384 11398 4386 11450
rect 4566 11398 4568 11450
rect 4322 11396 4328 11398
rect 4384 11396 4408 11398
rect 4464 11396 4488 11398
rect 4544 11396 4568 11398
rect 4624 11396 4630 11398
rect 4322 11387 4630 11396
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 4632 10606 4660 11086
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 3988 10198 4016 10542
rect 4252 10532 4304 10538
rect 4252 10474 4304 10480
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 4264 10130 4292 10474
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4322 10364 4630 10373
rect 4322 10362 4328 10364
rect 4384 10362 4408 10364
rect 4464 10362 4488 10364
rect 4544 10362 4568 10364
rect 4624 10362 4630 10364
rect 4384 10310 4386 10362
rect 4566 10310 4568 10362
rect 4322 10308 4328 10310
rect 4384 10308 4408 10310
rect 4464 10308 4488 10310
rect 4544 10308 4568 10310
rect 4624 10308 4630 10310
rect 4322 10299 4630 10308
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 4724 9722 4752 10406
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4816 9382 4844 10134
rect 4908 9586 4936 10542
rect 5092 10198 5120 11086
rect 5644 10606 5672 11222
rect 5736 11218 5764 12310
rect 6196 12170 6224 12650
rect 6380 12238 6408 12922
rect 6472 12866 6500 14418
rect 6564 12986 6592 15302
rect 7668 13938 7696 20046
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 7748 19780 7800 19786
rect 7748 19722 7800 19728
rect 7760 19378 7788 19722
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 8312 18970 8340 19790
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8392 18896 8444 18902
rect 8392 18838 8444 18844
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7760 18306 7788 18702
rect 7760 18290 8064 18306
rect 7760 18284 8076 18290
rect 7760 18278 8024 18284
rect 7760 18222 7788 18278
rect 8024 18226 8076 18232
rect 8404 18222 8432 18838
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8128 18086 8156 18158
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7760 15638 7788 16390
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 7748 15632 7800 15638
rect 7748 15574 7800 15580
rect 8128 15570 8156 15846
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6472 12838 6592 12866
rect 6564 12782 6592 12838
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6564 12434 6592 12718
rect 6564 12406 6776 12434
rect 6748 12306 6776 12406
rect 7024 12374 7052 13738
rect 7116 13734 7144 13806
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7116 13394 7144 13670
rect 8128 13462 8156 13874
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7116 12918 7144 13330
rect 7300 12986 7328 13330
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 8128 12850 8156 13398
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8404 12782 8432 13126
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 7116 12306 7144 12582
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 6380 12102 6408 12174
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 5828 11762 5856 12038
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6012 11218 6040 11630
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 4908 8566 4936 9522
rect 5000 9518 5028 9862
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5092 9110 5120 10134
rect 5184 9722 5212 10474
rect 5644 10130 5672 10542
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5276 9722 5304 10066
rect 5828 10062 5856 11154
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 5184 9058 5212 9318
rect 5276 9178 5304 9386
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5184 9030 5304 9058
rect 5368 9042 5396 9998
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 9518 5672 9862
rect 6012 9722 6040 11154
rect 6196 11150 6224 11222
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6196 10810 6224 11086
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6472 10606 6500 11562
rect 6656 11558 6684 11698
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6564 11218 6592 11494
rect 6748 11286 6776 12242
rect 7116 11898 7144 12242
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6840 11218 6868 11494
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6932 11014 6960 11766
rect 7116 11694 7144 11834
rect 7208 11694 7236 12378
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7392 11218 7420 12038
rect 7484 11762 7512 12106
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 7484 11354 7512 11698
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7668 11218 7696 11494
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 7116 10810 7144 11154
rect 8312 11150 8340 11698
rect 8404 11694 8432 12718
rect 8496 12714 8524 21286
rect 8588 20398 8616 21422
rect 9416 21078 9444 21626
rect 9600 21486 9628 22442
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9404 21072 9456 21078
rect 9404 21014 9456 21020
rect 9128 20800 9180 20806
rect 9128 20742 9180 20748
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 8680 20398 8708 20538
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 8576 19984 8628 19990
rect 8576 19926 8628 19932
rect 8588 17678 8616 19926
rect 8680 19310 8708 20334
rect 8944 20256 8996 20262
rect 8944 20198 8996 20204
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8956 18834 8984 20198
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8772 18426 8800 18702
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 8864 18222 8892 18770
rect 8956 18306 8984 18770
rect 8956 18278 9076 18306
rect 9048 18222 9076 18278
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8588 16726 8616 17614
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8864 17134 8892 17478
rect 9036 17264 9088 17270
rect 9036 17206 9088 17212
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8588 16046 8616 16662
rect 9048 16114 9076 17206
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 9048 15570 9076 16050
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 9140 14958 9168 20742
rect 9416 19310 9444 21014
rect 9692 21010 9720 21898
rect 9784 21486 9812 22442
rect 9864 22432 9916 22438
rect 9968 22386 9996 22646
rect 10428 22574 10456 22714
rect 10980 22642 11008 23054
rect 11072 22710 11100 23122
rect 11060 22704 11112 22710
rect 11112 22652 11192 22658
rect 11060 22646 11192 22652
rect 10968 22636 11020 22642
rect 11072 22630 11192 22646
rect 10968 22578 11020 22584
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 9916 22380 9996 22386
rect 9864 22374 9996 22380
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 9876 22358 9996 22374
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 9876 21622 9904 22034
rect 9864 21616 9916 21622
rect 9864 21558 9916 21564
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9784 21146 9812 21286
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9496 21004 9548 21010
rect 9496 20946 9548 20952
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9508 20806 9536 20946
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9692 20398 9720 20946
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9772 19916 9824 19922
rect 9876 19904 9904 21558
rect 9968 21010 9996 22358
rect 10060 22166 10088 22374
rect 10048 22160 10100 22166
rect 10048 22102 10100 22108
rect 10980 22030 11008 22578
rect 11060 22500 11112 22506
rect 11060 22442 11112 22448
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 10152 20602 10180 21898
rect 10244 21486 10272 21966
rect 10876 21616 10928 21622
rect 10876 21558 10928 21564
rect 10232 21480 10284 21486
rect 10232 21422 10284 21428
rect 10784 21480 10836 21486
rect 10784 21422 10836 21428
rect 10796 21350 10824 21422
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10796 21146 10824 21286
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 10336 20874 10364 20946
rect 10324 20868 10376 20874
rect 10324 20810 10376 20816
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 9824 19876 9904 19904
rect 9772 19858 9824 19864
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9416 18834 9444 19246
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9508 18766 9536 19722
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9324 16658 9352 17070
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9416 15094 9444 18566
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9508 16794 9536 17274
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9404 15088 9456 15094
rect 9404 15030 9456 15036
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9232 14482 9260 14962
rect 9416 14958 9444 15030
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9600 14482 9628 19110
rect 9784 18222 9812 19858
rect 10060 18902 10088 20334
rect 10336 19922 10364 20810
rect 10796 20602 10824 20946
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 10888 20466 10916 21558
rect 11072 21010 11100 22442
rect 11164 22098 11192 22630
rect 11256 22166 11284 23122
rect 11900 22574 11928 23122
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 13556 22642 13584 22918
rect 14292 22778 14320 22918
rect 14004 22772 14056 22778
rect 14004 22714 14056 22720
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 13912 22704 13964 22710
rect 13912 22646 13964 22652
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 11612 22568 11664 22574
rect 11348 22506 11560 22522
rect 11612 22510 11664 22516
rect 11888 22568 11940 22574
rect 11888 22510 11940 22516
rect 12072 22568 12124 22574
rect 12072 22510 12124 22516
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 11348 22500 11572 22506
rect 11348 22494 11520 22500
rect 11244 22160 11296 22166
rect 11244 22102 11296 22108
rect 11152 22092 11204 22098
rect 11152 22034 11204 22040
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 11164 20806 11192 22034
rect 11348 21962 11376 22494
rect 11520 22442 11572 22448
rect 11428 22432 11480 22438
rect 11428 22374 11480 22380
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11348 20806 11376 21898
rect 11440 21010 11468 22374
rect 11624 22234 11652 22510
rect 11612 22228 11664 22234
rect 11612 22170 11664 22176
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11624 20942 11652 22170
rect 11900 22166 11928 22510
rect 11888 22160 11940 22166
rect 11888 22102 11940 22108
rect 12084 22098 12112 22510
rect 11796 22092 11848 22098
rect 11716 22052 11796 22080
rect 11716 21146 11744 22052
rect 11796 22034 11848 22040
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 12070 21992 12126 22001
rect 12070 21927 12126 21936
rect 12084 21554 12112 21927
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 11704 21140 11756 21146
rect 11704 21082 11756 21088
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11336 20800 11388 20806
rect 11336 20742 11388 20748
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10980 19718 11008 20334
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10980 19310 11008 19654
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10048 18896 10100 18902
rect 10048 18838 10100 18844
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9692 17134 9720 17682
rect 9876 17270 9904 18022
rect 10060 17542 10088 18566
rect 10152 17678 10180 19110
rect 10980 18834 11008 19246
rect 11072 19242 11100 19858
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10336 18222 10364 18702
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10336 17882 10364 18158
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9692 16658 9720 17070
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9692 15570 9720 15982
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9784 15026 9812 16934
rect 9876 16726 9904 17206
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9968 16794 9996 16934
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 10060 16454 10088 17478
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10152 16266 10180 17614
rect 10244 17202 10272 17682
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10428 17134 10456 18362
rect 10612 18358 10640 18770
rect 10600 18352 10652 18358
rect 10968 18352 11020 18358
rect 10600 18294 10652 18300
rect 10888 18312 10968 18340
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10796 17134 10824 17750
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 9968 16238 10180 16266
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9784 14906 9812 14962
rect 9968 14958 9996 16238
rect 10140 15428 10192 15434
rect 10140 15370 10192 15376
rect 9692 14878 9812 14906
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 10152 14890 10180 15370
rect 10140 14884 10192 14890
rect 9692 14550 9720 14878
rect 10060 14844 10140 14872
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9048 13870 9076 14350
rect 9232 14006 9260 14418
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9416 13870 9444 14418
rect 9784 14414 9812 14758
rect 10060 14482 10088 14844
rect 10140 14826 10192 14832
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9048 13376 9076 13806
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9508 13462 9536 13670
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9600 13394 9628 14010
rect 9784 13870 9812 14350
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9968 13870 9996 14214
rect 10060 14006 10088 14418
rect 10152 14278 10180 14554
rect 10244 14482 10272 16390
rect 10784 16040 10836 16046
rect 10888 16028 10916 18312
rect 10968 18294 11020 18300
rect 11072 18154 11100 19178
rect 11256 18970 11284 19790
rect 11992 19310 12020 21490
rect 12176 21350 12204 21626
rect 12268 21554 12296 22510
rect 12808 22500 12860 22506
rect 12808 22442 12860 22448
rect 12820 22234 12848 22442
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 12716 22092 12768 22098
rect 12716 22034 12768 22040
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12636 21622 12664 21830
rect 12624 21616 12676 21622
rect 12624 21558 12676 21564
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12728 21418 12756 22034
rect 12820 21486 12848 22170
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12716 21412 12768 21418
rect 12716 21354 12768 21360
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12360 21146 12388 21354
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 12360 19854 12388 20402
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12452 19922 12480 20334
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 11980 19304 12032 19310
rect 11900 19252 11980 19258
rect 11900 19246 12032 19252
rect 11900 19230 12020 19246
rect 12348 19236 12400 19242
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11348 18426 11376 18770
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11336 18420 11388 18426
rect 11336 18362 11388 18368
rect 11624 18222 11652 18566
rect 11716 18358 11744 18770
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11900 18154 11928 19230
rect 12348 19178 12400 19184
rect 12072 18896 12124 18902
rect 12070 18864 12072 18873
rect 12124 18864 12126 18873
rect 12070 18799 12126 18808
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11992 18222 12020 18702
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 12084 17746 12112 18799
rect 12360 18222 12388 19178
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 10980 17338 11008 17682
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12360 17338 12388 17614
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12544 16046 12572 17682
rect 13004 16182 13032 21830
rect 13096 21690 13124 21966
rect 13084 21684 13136 21690
rect 13084 21626 13136 21632
rect 13188 21010 13216 22578
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 13280 21622 13308 22510
rect 13452 22500 13504 22506
rect 13452 22442 13504 22448
rect 13360 22432 13412 22438
rect 13360 22374 13412 22380
rect 13268 21616 13320 21622
rect 13268 21558 13320 21564
rect 13372 21486 13400 22374
rect 13464 22098 13492 22442
rect 13452 22092 13504 22098
rect 13452 22034 13504 22040
rect 13464 21690 13492 22034
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13556 21554 13584 22578
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 13648 21962 13676 22510
rect 13832 22030 13860 22578
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13636 21956 13688 21962
rect 13636 21898 13688 21904
rect 13728 21616 13780 21622
rect 13728 21558 13780 21564
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13360 21480 13412 21486
rect 13360 21422 13412 21428
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 13740 20806 13768 21558
rect 13924 21010 13952 22646
rect 14016 21486 14044 22714
rect 14476 22506 14504 23190
rect 16408 23186 16436 23600
rect 19536 23254 19564 23718
rect 22282 23600 22338 24000
rect 19708 23316 19760 23322
rect 19708 23258 19760 23264
rect 18144 23248 18196 23254
rect 18144 23190 18196 23196
rect 18696 23248 18748 23254
rect 18696 23190 18748 23196
rect 19524 23248 19576 23254
rect 19524 23190 19576 23196
rect 15108 23180 15160 23186
rect 15108 23122 15160 23128
rect 16396 23180 16448 23186
rect 16396 23122 16448 23128
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14464 22500 14516 22506
rect 14464 22442 14516 22448
rect 14660 22098 14688 22510
rect 15120 22506 15148 23122
rect 16028 23044 16080 23050
rect 16028 22986 16080 22992
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15108 22500 15160 22506
rect 15108 22442 15160 22448
rect 14924 22432 14976 22438
rect 14924 22374 14976 22380
rect 14936 22234 14964 22374
rect 14924 22228 14976 22234
rect 14924 22170 14976 22176
rect 14096 22092 14148 22098
rect 14096 22034 14148 22040
rect 14648 22092 14700 22098
rect 14648 22034 14700 22040
rect 14108 22001 14136 22034
rect 15016 22024 15068 22030
rect 14094 21992 14150 22001
rect 15016 21966 15068 21972
rect 14094 21927 14150 21936
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 14188 21344 14240 21350
rect 14188 21286 14240 21292
rect 14108 21146 14136 21286
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 13912 21004 13964 21010
rect 13912 20946 13964 20952
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 13188 19922 13216 20538
rect 14108 20466 14136 21082
rect 14200 20777 14228 21286
rect 14186 20768 14242 20777
rect 14186 20703 14242 20712
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13648 19990 13676 20198
rect 13636 19984 13688 19990
rect 13636 19926 13688 19932
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 13648 19446 13676 19926
rect 13740 19854 13768 20334
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13832 19922 13860 20198
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13832 19700 13860 19858
rect 13740 19672 13860 19700
rect 13636 19440 13688 19446
rect 13636 19382 13688 19388
rect 13648 18834 13676 19382
rect 13740 19310 13768 19672
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13820 19304 13872 19310
rect 13924 19292 13952 19858
rect 14108 19310 14136 19858
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14292 19310 14320 19790
rect 14384 19718 14412 20402
rect 14476 20398 14504 21422
rect 14660 20602 14688 21490
rect 14740 21480 14792 21486
rect 14738 21448 14740 21457
rect 14792 21448 14794 21457
rect 14738 21383 14794 21392
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 14844 19854 14872 21830
rect 14924 21072 14976 21078
rect 14924 21014 14976 21020
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14740 19780 14792 19786
rect 14740 19722 14792 19728
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14752 19310 14780 19722
rect 13872 19264 13952 19292
rect 14096 19304 14148 19310
rect 13820 19246 13872 19252
rect 14096 19246 14148 19252
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14556 19304 14608 19310
rect 14740 19304 14792 19310
rect 14556 19246 14608 19252
rect 14660 19264 14740 19292
rect 13740 18834 13768 19246
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13832 18698 13860 19246
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18970 14504 19110
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 13820 18692 13872 18698
rect 13820 18634 13872 18640
rect 14384 18358 14412 18770
rect 14464 18692 14516 18698
rect 14464 18634 14516 18640
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 13280 17678 13308 18294
rect 14476 17882 14504 18634
rect 14568 18426 14596 19246
rect 14660 18902 14688 19264
rect 14740 19246 14792 19252
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14648 18896 14700 18902
rect 14648 18838 14700 18844
rect 14752 18834 14780 19110
rect 14936 18952 14964 21014
rect 15028 21010 15056 21966
rect 15212 21962 15240 22714
rect 15752 22704 15804 22710
rect 15752 22646 15804 22652
rect 15764 22522 15792 22646
rect 16040 22642 16068 22986
rect 17500 22976 17552 22982
rect 17500 22918 17552 22924
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 16408 22574 16436 22714
rect 16764 22704 16816 22710
rect 16764 22646 16816 22652
rect 16856 22704 16908 22710
rect 16856 22646 16908 22652
rect 16396 22568 16448 22574
rect 15764 22494 16160 22522
rect 16396 22510 16448 22516
rect 15292 22432 15344 22438
rect 15752 22432 15804 22438
rect 15344 22409 15424 22420
rect 15344 22400 15438 22409
rect 15344 22392 15382 22400
rect 15292 22374 15344 22380
rect 15752 22374 15804 22380
rect 15382 22335 15438 22344
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 14844 18924 14964 18952
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 14844 17218 14872 18924
rect 15120 18834 15148 19654
rect 15108 18828 15160 18834
rect 14936 18788 15108 18816
rect 14936 18222 14964 18788
rect 15108 18770 15160 18776
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15108 18624 15160 18630
rect 15108 18566 15160 18572
rect 15028 18465 15056 18566
rect 15014 18456 15070 18465
rect 15014 18391 15070 18400
rect 15120 18306 15148 18566
rect 15028 18290 15148 18306
rect 15016 18284 15148 18290
rect 15068 18278 15148 18284
rect 15016 18226 15068 18232
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 15028 17338 15056 18226
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 14844 17190 15056 17218
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14464 17060 14516 17066
rect 14464 17002 14516 17008
rect 14476 16794 14504 17002
rect 14660 16998 14688 17070
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14464 16516 14516 16522
rect 14464 16458 14516 16464
rect 12992 16176 13044 16182
rect 12992 16118 13044 16124
rect 13004 16046 13032 16118
rect 14476 16046 14504 16458
rect 10836 16000 10916 16028
rect 12532 16040 12584 16046
rect 10784 15982 10836 15988
rect 12532 15982 12584 15988
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10336 15570 10364 15914
rect 10796 15706 10824 15982
rect 12256 15972 12308 15978
rect 12256 15914 12308 15920
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10428 15484 10456 15642
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 10692 15496 10744 15502
rect 10428 15456 10692 15484
rect 10692 15438 10744 15444
rect 11348 15366 11376 15574
rect 11992 15570 12020 15846
rect 12268 15706 12296 15914
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12268 15570 12296 15642
rect 12912 15570 12940 15846
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 11532 15366 11560 15506
rect 11900 15434 11928 15506
rect 11888 15428 11940 15434
rect 11888 15370 11940 15376
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10336 14362 10364 14894
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10244 14346 10364 14362
rect 10232 14340 10364 14346
rect 10284 14334 10364 14340
rect 10232 14282 10284 14288
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10152 13530 10180 13670
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10244 13394 10272 14282
rect 10612 13870 10640 14758
rect 10888 14482 10916 14758
rect 10980 14618 11008 15098
rect 11532 14958 11560 15302
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11336 14884 11388 14890
rect 11336 14826 11388 14832
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11348 14550 11376 14826
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10888 13954 10916 14214
rect 11348 14074 11376 14486
rect 11440 14414 11468 14758
rect 11624 14482 11652 15302
rect 11900 14906 11928 15370
rect 11992 15162 12020 15506
rect 12544 15162 12572 15506
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 11808 14878 11928 14906
rect 12728 14890 12756 15506
rect 12912 14890 12940 15506
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 12716 14884 12768 14890
rect 11808 14822 11836 14878
rect 12716 14826 12768 14832
rect 12900 14884 12952 14890
rect 12900 14826 12952 14832
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 11900 14618 11928 14758
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 12360 14482 12388 14758
rect 13096 14482 13124 15030
rect 13556 14958 13584 15302
rect 13832 15162 13860 15438
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 12348 14476 12400 14482
rect 13084 14476 13136 14482
rect 12348 14418 12400 14424
rect 13004 14436 13084 14464
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 10888 13926 11008 13954
rect 10980 13870 11008 13926
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 9220 13388 9272 13394
rect 9048 13348 9220 13376
rect 9220 13330 9272 13336
rect 9312 13388 9364 13394
rect 9588 13388 9640 13394
rect 9364 13348 9444 13376
rect 9312 13330 9364 13336
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8680 11694 8708 12718
rect 9048 12714 9076 13126
rect 9232 12714 9260 13330
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8956 12434 8984 12582
rect 8772 12406 8984 12434
rect 8772 11762 8800 12406
rect 9324 12238 9352 13194
rect 9416 12646 9444 13348
rect 9588 13330 9640 13336
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10152 12850 10180 13126
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 10244 12306 10272 13330
rect 10428 12782 10456 13670
rect 11808 13394 11836 14214
rect 12360 13938 12388 14282
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12360 13530 12388 13874
rect 13004 13870 13032 14436
rect 13084 14418 13136 14424
rect 13188 13938 13216 14554
rect 13452 14476 13504 14482
rect 13556 14464 13584 14894
rect 14108 14482 14136 14962
rect 14384 14958 14412 15846
rect 14660 15162 14688 16934
rect 15028 16658 15056 17190
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 14844 16250 14872 16594
rect 14922 16552 14978 16561
rect 14922 16487 14924 16496
rect 14976 16487 14978 16496
rect 14924 16458 14976 16464
rect 15028 16402 15056 16594
rect 14936 16374 15148 16402
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14936 16130 14964 16374
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 14844 16114 14964 16130
rect 14832 16108 14964 16114
rect 14884 16102 14964 16108
rect 14832 16050 14884 16056
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14752 15570 14780 15982
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14384 14618 14412 14894
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14660 14550 14688 14758
rect 15028 14618 15056 16186
rect 15120 16114 15148 16374
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15212 15094 15240 17002
rect 15304 15978 15332 21286
rect 15396 19174 15424 22335
rect 15568 22160 15620 22166
rect 15568 22102 15620 22108
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15488 21894 15516 21966
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 15488 21010 15516 21830
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15580 20534 15608 22102
rect 15764 22098 15792 22374
rect 16132 22098 16160 22494
rect 16408 22438 16436 22510
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16396 22432 16448 22438
rect 16500 22409 16528 22442
rect 16396 22374 16448 22380
rect 16486 22400 16542 22409
rect 16316 22234 16344 22374
rect 16486 22335 16542 22344
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16776 22098 16804 22646
rect 16868 22506 16896 22646
rect 17512 22506 17540 22918
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 17500 22500 17552 22506
rect 17500 22442 17552 22448
rect 17592 22500 17644 22506
rect 17592 22442 17644 22448
rect 17776 22500 17828 22506
rect 17776 22442 17828 22448
rect 17040 22160 17092 22166
rect 17040 22102 17092 22108
rect 15752 22092 15804 22098
rect 15752 22034 15804 22040
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16580 22092 16632 22098
rect 16580 22034 16632 22040
rect 16764 22092 16816 22098
rect 16764 22034 16816 22040
rect 15764 20942 15792 22034
rect 15936 21480 15988 21486
rect 15936 21422 15988 21428
rect 15948 21078 15976 21422
rect 16132 21418 16160 22034
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16120 21412 16172 21418
rect 16120 21354 16172 21360
rect 15936 21072 15988 21078
rect 15936 21014 15988 21020
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15948 20874 15976 21014
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 15936 20868 15988 20874
rect 15936 20810 15988 20816
rect 16316 20534 16344 20946
rect 15568 20528 15620 20534
rect 15568 20470 15620 20476
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16408 20466 16436 21422
rect 16500 21146 16528 21966
rect 16592 21457 16620 22034
rect 17052 21554 17080 22102
rect 17132 22092 17184 22098
rect 17132 22034 17184 22040
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17040 21548 17092 21554
rect 17040 21490 17092 21496
rect 17144 21486 17172 22034
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17132 21480 17184 21486
rect 16578 21448 16634 21457
rect 17132 21422 17184 21428
rect 16578 21383 16634 21392
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 17236 21010 17264 21626
rect 17420 21622 17448 22034
rect 17604 22030 17632 22442
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 17408 21616 17460 21622
rect 17408 21558 17460 21564
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17328 21146 17356 21422
rect 17420 21418 17448 21558
rect 17408 21412 17460 21418
rect 17408 21354 17460 21360
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17316 21140 17368 21146
rect 17316 21082 17368 21088
rect 17224 21004 17276 21010
rect 17224 20946 17276 20952
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 17512 20398 17540 21286
rect 17604 21010 17632 21966
rect 17788 21690 17816 22442
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17972 21894 18000 22374
rect 18156 22030 18184 23190
rect 18420 23180 18472 23186
rect 18420 23122 18472 23128
rect 18432 22506 18460 23122
rect 18708 22642 18736 23190
rect 19064 23180 19116 23186
rect 19064 23122 19116 23128
rect 18788 23112 18840 23118
rect 18788 23054 18840 23060
rect 18800 22710 18828 23054
rect 19076 22778 19104 23122
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 18788 22704 18840 22710
rect 18788 22646 18840 22652
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 19076 22522 19104 22714
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 18420 22500 18472 22506
rect 18420 22442 18472 22448
rect 18788 22500 18840 22506
rect 18788 22442 18840 22448
rect 18880 22500 18932 22506
rect 18880 22442 18932 22448
rect 18972 22500 19024 22506
rect 19076 22494 19196 22522
rect 18972 22442 19024 22448
rect 18800 22234 18828 22442
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17972 21486 18000 21830
rect 18248 21486 18276 22170
rect 18420 22160 18472 22166
rect 18420 22102 18472 22108
rect 18432 21554 18460 22102
rect 18892 21622 18920 22442
rect 18984 22098 19012 22442
rect 19064 22432 19116 22438
rect 19064 22374 19116 22380
rect 18972 22092 19024 22098
rect 18972 22034 19024 22040
rect 18880 21616 18932 21622
rect 18880 21558 18932 21564
rect 19076 21554 19104 22374
rect 19168 22098 19196 22494
rect 19156 22092 19208 22098
rect 19156 22034 19208 22040
rect 19260 22030 19288 22578
rect 19720 22098 19748 23258
rect 19892 23248 19944 23254
rect 19892 23190 19944 23196
rect 20076 23248 20128 23254
rect 20076 23190 20128 23196
rect 20996 23248 21048 23254
rect 20996 23190 21048 23196
rect 19904 23118 19932 23190
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 20088 22982 20116 23190
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 20076 22976 20128 22982
rect 20076 22918 20128 22924
rect 19996 22642 20024 22918
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 19800 22568 19852 22574
rect 19800 22510 19852 22516
rect 19812 22098 19840 22510
rect 20548 22506 20576 23054
rect 21008 22642 21036 23190
rect 22296 23186 22324 23600
rect 21088 23180 21140 23186
rect 21088 23122 21140 23128
rect 21364 23180 21416 23186
rect 21364 23122 21416 23128
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 21916 23180 21968 23186
rect 21916 23122 21968 23128
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 20536 22500 20588 22506
rect 20536 22442 20588 22448
rect 21008 22098 21036 22578
rect 19708 22092 19760 22098
rect 19708 22034 19760 22040
rect 19800 22092 19852 22098
rect 19800 22034 19852 22040
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19812 21894 19840 22034
rect 19800 21888 19852 21894
rect 19800 21830 19852 21836
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 19812 21690 19840 21830
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 18420 21548 18472 21554
rect 18420 21490 18472 21496
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 17960 21480 18012 21486
rect 17960 21422 18012 21428
rect 18236 21480 18288 21486
rect 18880 21480 18932 21486
rect 18236 21422 18288 21428
rect 18878 21448 18880 21457
rect 18932 21448 18934 21457
rect 18878 21383 18934 21392
rect 18892 21350 18920 21383
rect 18880 21344 18932 21350
rect 18880 21286 18932 21292
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 18328 20392 18380 20398
rect 18328 20334 18380 20340
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 17144 19922 17172 20198
rect 18156 20058 18184 20198
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15488 19242 15516 19314
rect 16408 19310 16436 19858
rect 18340 19786 18368 20334
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18432 19922 18460 19994
rect 18524 19922 18552 20198
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 18420 19916 18472 19922
rect 18420 19858 18472 19864
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18800 19854 18828 19994
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 17960 19780 18012 19786
rect 17960 19722 18012 19728
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 17972 19310 18000 19722
rect 18340 19446 18368 19722
rect 18892 19514 18920 20334
rect 19260 20058 19288 21490
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 21010 20484 21286
rect 20548 21010 20576 21422
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20536 21004 20588 21010
rect 20536 20946 20588 20952
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 20272 19922 20300 20742
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 19800 19916 19852 19922
rect 19800 19858 19852 19864
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 19064 19712 19116 19718
rect 19064 19654 19116 19660
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18880 19508 18932 19514
rect 18880 19450 18932 19456
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16396 19304 16448 19310
rect 16396 19246 16448 19252
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 15476 19236 15528 19242
rect 15476 19178 15528 19184
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 15396 18222 15424 18770
rect 15488 18737 15516 19178
rect 16316 18766 16344 19246
rect 16408 18902 16436 19246
rect 18236 19168 18288 19174
rect 18236 19110 18288 19116
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18248 18902 18276 19110
rect 16396 18896 16448 18902
rect 16394 18864 16396 18873
rect 18236 18896 18288 18902
rect 16448 18864 16450 18873
rect 18236 18838 18288 18844
rect 16394 18799 16450 18808
rect 18524 18766 18552 19110
rect 18708 18834 18736 19450
rect 19076 19310 19104 19654
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 16304 18760 16356 18766
rect 15474 18728 15530 18737
rect 16304 18702 16356 18708
rect 18512 18760 18564 18766
rect 18880 18760 18932 18766
rect 18564 18720 18644 18748
rect 18512 18702 18564 18708
rect 15474 18663 15530 18672
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 15384 17264 15436 17270
rect 15384 17206 15436 17212
rect 15396 16658 15424 17206
rect 15488 16810 15516 18090
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15580 17202 15608 18022
rect 15672 17746 15700 18158
rect 15764 17746 15792 18226
rect 16132 18222 16160 18634
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 16394 18456 16450 18465
rect 16394 18391 16450 18400
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 16040 17610 16068 17818
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16028 17604 16080 17610
rect 15856 17564 16028 17592
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15488 16782 15608 16810
rect 15476 16720 15528 16726
rect 15476 16662 15528 16668
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15488 16250 15516 16662
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15304 15638 15332 15914
rect 15292 15632 15344 15638
rect 15292 15574 15344 15580
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 14648 14544 14700 14550
rect 14648 14486 14700 14492
rect 13504 14436 13584 14464
rect 14096 14476 14148 14482
rect 13452 14418 13504 14424
rect 14096 14418 14148 14424
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 13084 13796 13136 13802
rect 13084 13738 13136 13744
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 11072 12434 11100 12922
rect 11152 12436 11204 12442
rect 11072 12406 11152 12434
rect 11152 12378 11204 12384
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8404 11150 8432 11630
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8588 11286 8616 11494
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8312 11014 8340 11086
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 8312 10674 8340 10950
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8404 10606 8432 11086
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 6368 10532 6420 10538
rect 6368 10474 6420 10480
rect 6380 10266 6408 10474
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6472 9926 6500 10542
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6748 9722 6776 10406
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6932 9722 6960 10066
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6932 9110 6960 9386
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7576 9178 7604 9318
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 7668 9092 7696 9454
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 7748 9104 7800 9110
rect 7668 9064 7748 9092
rect 5276 8974 5304 9030
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 4448 7546 4476 7958
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4540 7342 4568 7890
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4264 7002 4292 7278
rect 4724 7274 4752 8230
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 5000 7546 5028 7754
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 5092 7274 5120 7822
rect 5276 7818 5304 8910
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 4724 6458 4752 7210
rect 5184 6934 5212 7686
rect 5368 7342 5396 8978
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 8634 7144 8774
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7668 8430 7696 9064
rect 7748 9046 7800 9052
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7852 8634 7880 9046
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 5644 7886 5672 8366
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 5276 6662 5304 7278
rect 5644 7002 5672 7822
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5920 6866 5948 8026
rect 6012 7970 6040 8230
rect 6012 7942 6132 7970
rect 6932 7954 6960 8230
rect 6104 7886 6132 7942
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6288 7546 6316 7822
rect 6840 7750 6868 7890
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6840 7478 6868 7686
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6840 6934 6868 7414
rect 6932 7274 6960 7754
rect 7116 7342 7144 7890
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6932 7002 6960 7210
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 7116 6866 7144 7278
rect 7484 7274 7512 8298
rect 7852 8090 7880 8570
rect 8220 8090 8248 9318
rect 8404 8634 8432 9454
rect 8588 9450 8616 11222
rect 8680 10130 8708 11630
rect 8772 11082 8800 11698
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8588 8906 8616 9386
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8220 7546 8248 8026
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8312 7342 8340 8502
rect 8484 8424 8536 8430
rect 8588 8412 8616 8842
rect 8680 8838 8708 10066
rect 8772 9110 8800 10066
rect 8864 10062 8892 10610
rect 9232 10470 9260 11494
rect 9416 11354 9444 11562
rect 9876 11354 9904 12038
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9324 10198 9352 11290
rect 10244 11218 10272 11630
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10336 11150 10364 11494
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 10810 9536 10950
rect 9496 10804 9548 10810
rect 9956 10804 10008 10810
rect 9496 10746 9548 10752
rect 9784 10764 9956 10792
rect 9784 10606 9812 10764
rect 9956 10746 10008 10752
rect 10336 10606 10364 11086
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9692 10130 9720 10406
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 9784 9518 9812 10542
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8430 8708 8774
rect 8536 8384 8616 8412
rect 8668 8424 8720 8430
rect 8484 8366 8536 8372
rect 8668 8366 8720 8372
rect 8680 7954 8708 8366
rect 8956 8022 8984 9318
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9324 8090 9352 8298
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 8944 8016 8996 8022
rect 8944 7958 8996 7964
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8680 7478 8708 7890
rect 9508 7750 9536 9318
rect 9784 9178 9812 9454
rect 9968 9178 9996 9658
rect 10336 9586 10364 10406
rect 10428 9926 10456 10678
rect 10520 10606 10548 10746
rect 11072 10606 11100 11086
rect 11164 11014 11192 12378
rect 11624 12374 11652 13126
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11348 11626 11376 12174
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 11256 11354 11284 11562
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9600 8906 9628 8978
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9784 8634 9812 9114
rect 10796 9042 10824 9114
rect 10888 9042 10916 9386
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10152 8022 10180 8298
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5828 6458 5856 6734
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 7392 6186 7420 7142
rect 7760 7002 7788 7210
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 8680 6322 8708 7414
rect 10152 6934 10180 7958
rect 10140 6928 10192 6934
rect 10140 6870 10192 6876
rect 10244 6662 10272 8774
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10336 8090 10364 8570
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10428 7002 10456 7142
rect 10612 7002 10640 8774
rect 10704 8498 10732 8842
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10796 7954 10824 8978
rect 10888 8022 10916 8978
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 11072 8022 11100 8502
rect 11256 8498 11284 8774
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11348 8430 11376 11562
rect 11716 11354 11744 12582
rect 11992 12442 12020 13262
rect 12084 12986 12112 13262
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12348 12776 12400 12782
rect 12452 12764 12480 13466
rect 12820 13394 12848 13670
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12400 12736 12480 12764
rect 12348 12718 12400 12724
rect 12544 12646 12572 13262
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12782 12756 13126
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12636 12442 12664 12650
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 12360 11150 12388 11494
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11532 10606 11560 10950
rect 12360 10606 12388 11086
rect 12544 10810 12572 11154
rect 12636 11014 12664 12378
rect 12728 11218 12756 12582
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12636 10742 12664 10950
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12728 10606 12756 11154
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 11624 10062 11652 10406
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11612 9036 11664 9042
rect 11716 9024 11744 10066
rect 12176 9586 12204 10406
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12268 9722 12296 9998
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12452 9654 12480 10066
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 12084 9178 12112 9454
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11664 8996 11744 9024
rect 12808 9036 12860 9042
rect 11612 8978 11664 8984
rect 12808 8978 12860 8984
rect 11624 8906 11652 8978
rect 11612 8900 11664 8906
rect 11612 8842 11664 8848
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11348 8022 11376 8366
rect 11624 8090 11652 8842
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8634 12480 8774
rect 12820 8634 12848 8978
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 13004 8362 13032 9318
rect 13096 9110 13124 13738
rect 13280 13530 13308 13874
rect 13740 13870 13768 14214
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13740 13394 13768 13806
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13372 12306 13400 12718
rect 13832 12306 13860 13942
rect 14108 13870 14136 14418
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14108 13394 14136 13670
rect 14096 13388 14148 13394
rect 14292 13376 14320 14214
rect 14384 13870 14412 14214
rect 14660 14074 14688 14214
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14372 13388 14424 13394
rect 14292 13348 14372 13376
rect 14096 13330 14148 13336
rect 14372 13330 14424 13336
rect 14832 13388 14884 13394
rect 14936 13376 14964 13874
rect 15488 13870 15516 14894
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 14884 13348 14964 13376
rect 14832 13330 14884 13336
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13924 12306 13952 13262
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14200 12782 14228 13126
rect 14936 12918 14964 13348
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15304 12986 15332 13262
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 14924 12912 14976 12918
rect 14924 12854 14976 12860
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 15304 12434 15332 12922
rect 15488 12714 15516 13806
rect 15580 12850 15608 16782
rect 15856 16590 15884 17564
rect 16028 17546 16080 17552
rect 16132 17134 16160 17750
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16132 16658 16160 17070
rect 16224 16998 16252 17478
rect 16316 17202 16344 17614
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16120 16652 16172 16658
rect 16040 16612 16120 16640
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15936 16584 15988 16590
rect 16040 16572 16068 16612
rect 16120 16594 16172 16600
rect 15988 16544 16068 16572
rect 15936 16526 15988 16532
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16132 16046 16160 16390
rect 16224 16046 16252 16662
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16132 14958 16160 15438
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 16132 13530 16160 13738
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16408 13326 16436 18391
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16500 17270 16528 17614
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16776 17134 16804 18022
rect 16868 17746 16896 18022
rect 17132 17808 17184 17814
rect 17132 17750 17184 17756
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 17144 17338 17172 17750
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 16948 17264 17000 17270
rect 16948 17206 17000 17212
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16684 16794 16712 17070
rect 16868 17066 16896 17138
rect 16856 17060 16908 17066
rect 16856 17002 16908 17008
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16776 16658 16804 16934
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16488 16040 16540 16046
rect 16592 16028 16620 16458
rect 16684 16250 16712 16594
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 16540 16000 16620 16028
rect 16488 15982 16540 15988
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16500 13258 16528 15982
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16684 15638 16712 15846
rect 16672 15632 16724 15638
rect 16672 15574 16724 15580
rect 16776 14958 16804 15846
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16592 13734 16620 14418
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 13870 16804 14214
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16592 13462 16620 13670
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15212 12406 15332 12434
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14108 11694 14136 12174
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 14832 12096 14884 12102
rect 15120 12050 15148 12106
rect 14832 12038 14884 12044
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13740 11082 13768 11154
rect 14844 11082 14872 12038
rect 15028 12022 15148 12050
rect 15028 11626 15056 12022
rect 15212 11626 15240 12406
rect 15396 11694 15424 12582
rect 15764 11898 15792 12582
rect 16592 12374 16620 13398
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16776 12238 16804 13806
rect 16868 13326 16896 16186
rect 16960 16046 16988 17206
rect 17144 17066 17172 17274
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17144 16658 17172 17002
rect 17328 16726 17356 17614
rect 17420 17338 17448 17682
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17512 17202 17540 18158
rect 17592 18148 17644 18154
rect 17592 18090 17644 18096
rect 17604 17610 17632 18090
rect 17696 17882 17724 18158
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17604 17134 17632 17546
rect 17696 17338 17724 17818
rect 18524 17814 18552 18566
rect 18616 18358 18644 18720
rect 18880 18702 18932 18708
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18708 18290 18736 18566
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18800 18222 18828 18566
rect 18892 18222 18920 18702
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18512 17808 18564 17814
rect 18512 17750 18564 17756
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 18064 17202 18092 17478
rect 18156 17338 18184 17614
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17328 16590 17356 16662
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17052 16046 17080 16390
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 17420 15570 17448 17002
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16250 17540 16934
rect 18248 16794 18276 17682
rect 18328 17604 18380 17610
rect 18328 17546 18380 17552
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18340 16522 18368 17546
rect 18616 17134 18644 18158
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18708 17746 18736 18022
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18696 17604 18748 17610
rect 18696 17546 18748 17552
rect 18708 17134 18736 17546
rect 18984 17338 19012 18226
rect 19352 18222 19380 19178
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18432 16658 18460 17070
rect 18616 16658 18644 17070
rect 19352 16998 19380 18158
rect 19536 17746 19564 18702
rect 19812 18426 19840 19858
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20272 19446 20300 19654
rect 20260 19440 20312 19446
rect 20260 19382 20312 19388
rect 20260 19304 20312 19310
rect 20364 19292 20392 19994
rect 20456 19446 20484 20198
rect 20548 19802 20576 20334
rect 20640 19922 20668 21830
rect 21008 21486 21036 22034
rect 21100 21486 21128 23122
rect 21376 22982 21404 23122
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 21088 21480 21140 21486
rect 21088 21422 21140 21428
rect 20732 21010 20760 21422
rect 21008 21078 21036 21422
rect 21192 21418 21220 21898
rect 21376 21486 21404 22918
rect 21468 22778 21496 23122
rect 21732 22976 21784 22982
rect 21732 22918 21784 22924
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21548 22432 21600 22438
rect 21548 22374 21600 22380
rect 21640 22432 21692 22438
rect 21640 22374 21692 22380
rect 21560 22234 21588 22374
rect 21548 22228 21600 22234
rect 21548 22170 21600 22176
rect 21456 22160 21508 22166
rect 21456 22102 21508 22108
rect 21468 21690 21496 22102
rect 21560 22098 21588 22170
rect 21652 22098 21680 22374
rect 21548 22092 21600 22098
rect 21548 22034 21600 22040
rect 21640 22092 21692 22098
rect 21640 22034 21692 22040
rect 21744 22012 21772 22918
rect 21928 22778 21956 23122
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 22008 22704 22060 22710
rect 22008 22646 22060 22652
rect 21824 22024 21876 22030
rect 21744 21984 21824 22012
rect 21744 21978 21772 21984
rect 21560 21962 21772 21978
rect 21824 21966 21876 21972
rect 21548 21956 21772 21962
rect 21600 21950 21772 21956
rect 21548 21898 21600 21904
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21180 21412 21232 21418
rect 21180 21354 21232 21360
rect 20996 21072 21048 21078
rect 20996 21014 21048 21020
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20732 20058 20760 20334
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 21008 19854 21036 21014
rect 21744 21010 21772 21830
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 21100 20330 21128 20946
rect 21548 20936 21600 20942
rect 21836 20890 21864 21966
rect 21916 21956 21968 21962
rect 21916 21898 21968 21904
rect 21928 21418 21956 21898
rect 21916 21412 21968 21418
rect 21916 21354 21968 21360
rect 22020 21350 22048 22646
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22204 22030 22232 22442
rect 22572 22166 22600 22918
rect 22560 22160 22612 22166
rect 22560 22102 22612 22108
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 21548 20878 21600 20884
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 21088 20324 21140 20330
rect 21088 20266 21140 20272
rect 21284 20058 21312 20742
rect 21560 20602 21588 20878
rect 21744 20862 21864 20890
rect 22112 20874 22140 21830
rect 22204 21690 22232 21966
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22100 20868 22152 20874
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21468 20058 21496 20198
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 20996 19848 21048 19854
rect 20548 19786 20668 19802
rect 20996 19790 21048 19796
rect 20548 19780 20680 19786
rect 20548 19774 20628 19780
rect 20628 19722 20680 19728
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20640 19310 20668 19722
rect 21100 19310 21128 19858
rect 20312 19264 20392 19292
rect 20444 19304 20496 19310
rect 20260 19246 20312 19252
rect 20444 19246 20496 19252
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 19996 18902 20024 19110
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 19800 18420 19852 18426
rect 19800 18362 19852 18368
rect 19524 17740 19576 17746
rect 19524 17682 19576 17688
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16794 19380 16934
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18328 16516 18380 16522
rect 18328 16458 18380 16464
rect 19444 16250 19472 17478
rect 19536 17134 19564 17682
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19984 17060 20036 17066
rect 19984 17002 20036 17008
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19444 16114 19472 16186
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 18880 16040 18932 16046
rect 18880 15982 18932 15988
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17512 15706 17540 15914
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16960 14074 16988 14350
rect 17420 14278 17448 14418
rect 17512 14414 17540 15642
rect 17696 15570 17724 15982
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17696 15162 17724 15506
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17604 14550 17632 14758
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17684 14476 17736 14482
rect 17788 14464 17816 15302
rect 17880 14890 17908 15506
rect 18892 15502 18920 15982
rect 19536 15570 19564 15982
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19720 15570 19748 15846
rect 19904 15570 19932 15846
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19708 15564 19760 15570
rect 19708 15506 19760 15512
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17736 14436 17816 14464
rect 17684 14418 17736 14424
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17420 13462 17448 14214
rect 17880 14074 17908 14826
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17972 14074 18000 14418
rect 18432 14414 18460 15302
rect 18892 15162 18920 15438
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18708 14618 18736 14826
rect 18892 14618 18920 14826
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18064 14074 18092 14350
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17880 13818 17908 14010
rect 18156 13938 18184 14350
rect 18328 14340 18380 14346
rect 18328 14282 18380 14288
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 18340 13870 18368 14282
rect 18328 13864 18380 13870
rect 17592 13796 17644 13802
rect 17880 13790 18000 13818
rect 18328 13806 18380 13812
rect 17592 13738 17644 13744
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16868 12850 16896 13262
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16132 11898 16160 12038
rect 16592 11898 16620 12174
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 15752 11892 15804 11898
rect 15580 11852 15752 11880
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 13740 10606 13768 11018
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14568 10674 14596 10950
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14844 10606 14872 11018
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14936 10606 14964 10950
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14740 10532 14792 10538
rect 14740 10474 14792 10480
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10062 13768 10406
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 14556 10124 14608 10130
rect 14608 10084 14688 10112
rect 14556 10066 14608 10072
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13832 9450 13860 10066
rect 14660 9722 14688 10084
rect 14752 10062 14780 10474
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 13084 9104 13136 9110
rect 13832 9058 13860 9386
rect 13084 9046 13136 9052
rect 12992 8356 13044 8362
rect 12992 8298 13044 8304
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10888 7546 10916 7958
rect 10968 7880 11020 7886
rect 11348 7834 11376 7958
rect 13096 7954 13124 9046
rect 13740 9042 13860 9058
rect 14292 9042 14320 9386
rect 14476 9042 14504 9590
rect 14660 9330 14688 9658
rect 14752 9518 14780 9862
rect 14844 9722 14872 9862
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14660 9302 14780 9330
rect 14752 9042 14780 9302
rect 14936 9042 14964 9386
rect 15028 9042 15056 11562
rect 15212 11218 15240 11562
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15304 11218 15332 11494
rect 15580 11218 15608 11852
rect 15752 11834 15804 11840
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15120 10062 15148 10406
rect 16408 10266 16436 11222
rect 16592 11150 16620 11834
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16592 11014 16620 11086
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16684 10690 16712 11562
rect 16776 11354 16804 11834
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16868 11150 16896 12038
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16592 10662 16712 10690
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15212 9586 15240 9930
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15304 9518 15332 9862
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15396 9110 15424 10066
rect 16316 9518 16344 10066
rect 16408 9586 16436 10202
rect 16592 9654 16620 10662
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 16684 9654 16712 10474
rect 17052 10266 17080 11154
rect 17236 11082 17264 11630
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17224 11076 17276 11082
rect 17224 11018 17276 11024
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16776 9722 16804 9862
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16396 9580 16448 9586
rect 17040 9580 17092 9586
rect 16396 9522 16448 9528
rect 16776 9540 17040 9568
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 13728 9036 13860 9042
rect 13780 9030 13860 9036
rect 13728 8978 13780 8984
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13464 8362 13492 8774
rect 13832 8514 13860 9030
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 13740 8486 13860 8514
rect 13740 8430 13768 8486
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13372 8022 13400 8230
rect 13832 8090 13860 8486
rect 13924 8430 13952 8774
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 11020 7828 11376 7834
rect 10968 7822 11376 7828
rect 10980 7806 11376 7822
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 11072 7342 11100 7806
rect 14108 7546 14136 8774
rect 14752 8294 14780 8978
rect 14936 8362 14964 8978
rect 15028 8634 15056 8978
rect 15396 8974 15424 9046
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15028 8430 15056 8570
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14292 7342 14320 8230
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14476 7342 14504 8026
rect 14936 7342 14964 8298
rect 15120 7954 15148 8842
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15212 8090 15240 8774
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15304 7750 15332 8774
rect 15396 8634 15424 8910
rect 15488 8906 15516 9454
rect 16408 8906 16436 9522
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16408 8634 16436 8842
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 15476 8356 15528 8362
rect 16500 8344 16528 9454
rect 16776 9382 16804 9540
rect 17040 9522 17092 9528
rect 17328 9382 17356 11494
rect 17420 11354 17448 11630
rect 17604 11354 17632 13738
rect 17972 13734 18000 13790
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 17880 12782 17908 13398
rect 18156 12850 18184 13466
rect 18616 13190 18644 14418
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18984 13870 19012 14214
rect 19076 14074 19104 14758
rect 19260 14278 19288 15098
rect 19812 15026 19840 15302
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19352 14006 19380 14214
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19904 13870 19932 14894
rect 19996 13938 20024 17002
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20088 16726 20116 16934
rect 20076 16720 20128 16726
rect 20076 16662 20128 16668
rect 20088 16046 20116 16662
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17880 12442 17908 12718
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17972 12374 18000 12582
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17972 11626 18000 12038
rect 18064 11898 18092 12650
rect 18156 12374 18184 12786
rect 18616 12782 18644 13126
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 18156 11354 18184 12310
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 18248 11898 18276 12242
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18432 11626 18460 12582
rect 18616 12442 18644 12718
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18800 11830 18828 13806
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 19260 12714 19288 13398
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19352 12918 19380 13194
rect 19904 13190 19932 13670
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19720 12782 19748 13126
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 19248 12708 19300 12714
rect 19432 12708 19484 12714
rect 19300 12668 19380 12696
rect 19248 12650 19300 12656
rect 19076 12102 19104 12650
rect 19156 12640 19208 12646
rect 19208 12588 19288 12594
rect 19156 12582 19288 12588
rect 19168 12566 19288 12582
rect 19260 12434 19288 12566
rect 19168 12406 19288 12434
rect 19168 12238 19196 12406
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 18788 11824 18840 11830
rect 18788 11766 18840 11772
rect 18420 11620 18472 11626
rect 18420 11562 18472 11568
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 17604 10826 17632 11290
rect 18432 11286 18460 11562
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17512 10798 17632 10826
rect 17512 10742 17540 10798
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17512 9654 17540 10066
rect 17788 9722 17816 10202
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17880 9450 17908 11154
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18248 10606 18276 10950
rect 18340 10810 18368 10950
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 18156 10130 18184 10474
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 16868 8634 16896 9318
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16580 8356 16632 8362
rect 16500 8316 16580 8344
rect 15476 8298 15528 8304
rect 16580 8298 16632 8304
rect 17224 8356 17276 8362
rect 17328 8344 17356 9318
rect 18156 9110 18184 10066
rect 18432 9722 18460 11222
rect 19168 10606 19196 12174
rect 19352 11626 19380 12668
rect 19432 12650 19484 12656
rect 19444 11694 19472 12650
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19444 11354 19472 11494
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 19248 9716 19300 9722
rect 19248 9658 19300 9664
rect 18248 9110 18276 9658
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 18800 9178 18828 9318
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 18236 9104 18288 9110
rect 18236 9046 18288 9052
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17604 8634 17632 8978
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18340 8634 18368 8774
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 17276 8316 17356 8344
rect 17224 8298 17276 8304
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15396 8090 15424 8230
rect 15488 8090 15516 8298
rect 18432 8090 18460 8774
rect 18892 8498 18920 8774
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 19168 8430 19196 9318
rect 19260 9042 19288 9658
rect 19628 9518 19656 9862
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 19628 8022 19656 9454
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19720 8090 19748 9318
rect 19812 8906 19840 9318
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 19616 8016 19668 8022
rect 19616 7958 19668 7964
rect 19812 7954 19840 8842
rect 19904 8566 19932 9998
rect 19996 9382 20024 13874
rect 20180 13394 20208 19110
rect 20456 18426 20484 19246
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20548 18222 20576 18906
rect 21284 18902 21312 19110
rect 21272 18896 21324 18902
rect 21272 18838 21324 18844
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 20916 18290 20944 18566
rect 21560 18306 21588 18566
rect 21652 18426 21680 20266
rect 21744 19854 21772 20862
rect 22100 20810 22152 20816
rect 21916 20800 21968 20806
rect 21916 20742 21968 20748
rect 21928 20398 21956 20742
rect 22652 20528 22704 20534
rect 22652 20470 22704 20476
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 22192 20392 22244 20398
rect 22192 20334 22244 20340
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21744 19242 21772 19790
rect 21732 19236 21784 19242
rect 21732 19178 21784 19184
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 20904 18284 20956 18290
rect 21560 18278 21680 18306
rect 20904 18226 20956 18232
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20548 16658 20576 18158
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20364 15910 20392 16186
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20364 15366 20392 15846
rect 20456 15706 20484 15846
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20364 14890 20392 15302
rect 20456 14958 20484 15642
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20444 14952 20496 14958
rect 20444 14894 20496 14900
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 20548 14074 20576 15506
rect 20628 15496 20680 15502
rect 20680 15456 20760 15484
rect 20628 15438 20680 15444
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20640 15162 20668 15302
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20732 15026 20760 15456
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20824 14278 20852 17614
rect 20916 16046 20944 18226
rect 21652 18222 21680 18278
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 21284 17746 21312 18158
rect 21548 18148 21600 18154
rect 21548 18090 21600 18096
rect 21560 17882 21588 18090
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21272 17740 21324 17746
rect 21272 17682 21324 17688
rect 21652 17134 21680 18158
rect 21928 18086 21956 18770
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21928 17746 21956 18022
rect 21824 17740 21876 17746
rect 21824 17682 21876 17688
rect 21916 17740 21968 17746
rect 21916 17682 21968 17688
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 21284 16794 21312 17002
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 21744 16658 21772 16934
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21744 16182 21772 16594
rect 21732 16176 21784 16182
rect 21732 16118 21784 16124
rect 21744 16046 21772 16118
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21456 15972 21508 15978
rect 21456 15914 21508 15920
rect 20904 15632 20956 15638
rect 20904 15574 20956 15580
rect 20916 14890 20944 15574
rect 21468 15502 21496 15914
rect 21744 15570 21772 15982
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21284 15026 21312 15302
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 20904 14884 20956 14890
rect 20904 14826 20956 14832
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 20272 13190 20300 13806
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20548 13326 20576 13670
rect 20916 13546 20944 14826
rect 21468 14074 21496 14894
rect 21836 14618 21864 17682
rect 22204 17678 22232 20334
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22388 19922 22416 20198
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22296 19174 22324 19858
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 22112 17338 22140 17546
rect 22204 17338 22232 17614
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 22112 15502 22140 15914
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 22020 14958 22048 15370
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 20640 13518 20944 13546
rect 20640 13326 20668 13518
rect 20916 13462 20944 13518
rect 20720 13456 20772 13462
rect 20720 13398 20772 13404
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20548 12986 20576 13262
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20732 12442 20760 13398
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20824 13190 20852 13262
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20364 11354 20392 11834
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20732 11218 20760 12378
rect 20824 12306 20852 13126
rect 21100 12986 21128 13806
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21008 12306 21036 12922
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20168 9444 20220 9450
rect 20168 9386 20220 9392
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 8634 20024 9318
rect 20180 9178 20208 9386
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20076 9104 20128 9110
rect 20076 9046 20128 9052
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19892 8560 19944 8566
rect 20088 8537 20116 9046
rect 20272 9042 20300 10066
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20548 9110 20576 9318
rect 20444 9104 20496 9110
rect 20444 9046 20496 9052
rect 20536 9104 20588 9110
rect 20536 9046 20588 9052
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 20180 8838 20208 8978
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20456 8634 20484 9046
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 19892 8502 19944 8508
rect 20074 8528 20130 8537
rect 19904 8401 19932 8502
rect 20074 8463 20130 8472
rect 19890 8392 19946 8401
rect 19890 8327 19946 8336
rect 19904 8022 19932 8327
rect 20640 8090 20668 8978
rect 20732 8838 20760 10746
rect 21100 10690 21128 12242
rect 21192 11898 21220 13398
rect 21468 13190 21496 14010
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21284 12986 21312 13126
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21192 11150 21220 11834
rect 21284 11626 21312 12174
rect 21376 11694 21404 12718
rect 21456 12708 21508 12714
rect 21456 12650 21508 12656
rect 21468 12102 21496 12650
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21560 11778 21588 14418
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21652 13190 21680 13330
rect 21836 13326 21864 14554
rect 22112 14550 22140 15438
rect 22100 14544 22152 14550
rect 22100 14486 22152 14492
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 21928 14074 21956 14350
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 22112 13870 22140 14486
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 13462 22140 13670
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 22204 13326 22232 17070
rect 22296 16250 22324 19110
rect 22388 18970 22416 19858
rect 22664 19718 22692 20470
rect 22468 19712 22520 19718
rect 22468 19654 22520 19660
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22744 19712 22796 19718
rect 22744 19654 22796 19660
rect 23018 19680 23074 19689
rect 22480 19310 22508 19654
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 22572 18970 22600 19450
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22572 18170 22600 18906
rect 22572 18142 22692 18170
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22388 17746 22416 18022
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22296 14498 22324 15982
rect 22572 15910 22600 17682
rect 22664 16046 22692 18142
rect 22756 16726 22784 19654
rect 23018 19615 23074 19624
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22848 17678 22876 19246
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 22940 18086 22968 18770
rect 22928 18080 22980 18086
rect 22928 18022 22980 18028
rect 23032 17814 23060 19615
rect 23020 17808 23072 17814
rect 23020 17750 23072 17756
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 22744 16720 22796 16726
rect 22744 16662 22796 16668
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22664 15570 22692 15982
rect 22836 15904 22888 15910
rect 22836 15846 22888 15852
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22388 14958 22416 15302
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22560 14884 22612 14890
rect 22560 14826 22612 14832
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22296 14482 22416 14498
rect 22296 14476 22428 14482
rect 22296 14470 22376 14476
rect 22296 13870 22324 14470
rect 22376 14418 22428 14424
rect 22480 14346 22508 14758
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 21652 12782 21680 13126
rect 21640 12776 21692 12782
rect 21640 12718 21692 12724
rect 21732 12640 21784 12646
rect 21732 12582 21784 12588
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 21744 12374 21772 12582
rect 21732 12368 21784 12374
rect 21732 12310 21784 12316
rect 21928 12102 21956 12582
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21468 11750 21588 11778
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21272 11620 21324 11626
rect 21272 11562 21324 11568
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 21008 10662 21128 10690
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20824 9722 20852 10066
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20824 8566 20852 9658
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20732 8022 20760 8298
rect 19892 8016 19944 8022
rect 19892 7958 19944 7964
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 20824 7750 20852 8502
rect 20916 8294 20944 10066
rect 21008 9654 21036 10662
rect 21284 10554 21312 11562
rect 21088 10532 21140 10538
rect 21088 10474 21140 10480
rect 21192 10526 21312 10554
rect 21100 10198 21128 10474
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 20996 9648 21048 9654
rect 20996 9590 21048 9596
rect 21192 9518 21220 10526
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 21192 8974 21220 9454
rect 21284 9110 21312 10406
rect 21468 10266 21496 11750
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21560 11354 21588 11562
rect 21652 11354 21680 12038
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 22112 11218 22140 13126
rect 22204 12918 22232 13262
rect 22376 13252 22428 13258
rect 22572 13240 22600 14826
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 22428 13212 22600 13240
rect 22652 13252 22704 13258
rect 22376 13194 22428 13200
rect 22652 13194 22704 13200
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22296 11898 22324 12718
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22296 11286 22324 11834
rect 22388 11558 22416 13194
rect 22664 12306 22692 13194
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22376 11552 22428 11558
rect 22376 11494 22428 11500
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22388 11218 22416 11494
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 21456 10260 21508 10266
rect 21456 10202 21508 10208
rect 21548 10056 21600 10062
rect 21548 9998 21600 10004
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 21008 8430 21036 8774
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20916 8022 20944 8230
rect 20904 8016 20956 8022
rect 20904 7958 20956 7964
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20916 7342 20944 7958
rect 21192 7546 21220 8366
rect 21376 7954 21404 8910
rect 21560 8838 21588 9998
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 21836 9518 21864 9862
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21468 8294 21496 8434
rect 21560 8362 21588 8774
rect 21928 8566 21956 10542
rect 22020 10266 22048 10746
rect 22112 10606 22140 11154
rect 22756 10810 22784 14418
rect 22848 14346 22876 15846
rect 22928 14544 22980 14550
rect 22928 14486 22980 14492
rect 22836 14340 22888 14346
rect 22836 14282 22888 14288
rect 22744 10804 22796 10810
rect 22744 10746 22796 10752
rect 22560 10736 22612 10742
rect 22560 10678 22612 10684
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22008 10260 22060 10266
rect 22112 10248 22140 10542
rect 22192 10260 22244 10266
rect 22112 10220 22192 10248
rect 22008 10202 22060 10208
rect 22192 10202 22244 10208
rect 21916 8560 21968 8566
rect 21916 8502 21968 8508
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21548 8356 21600 8362
rect 21548 8298 21600 8304
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21652 8022 21680 8434
rect 21836 8401 21864 8434
rect 21822 8392 21878 8401
rect 21822 8327 21878 8336
rect 21928 8090 21956 8502
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 22020 8090 22048 8366
rect 22204 8362 22232 10202
rect 22388 8634 22416 10542
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22480 10130 22508 10406
rect 22468 10124 22520 10130
rect 22468 10066 22520 10072
rect 22572 9178 22600 10678
rect 22652 10600 22704 10606
rect 22652 10542 22704 10548
rect 22664 10130 22692 10542
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22664 9382 22692 10066
rect 22848 9994 22876 14282
rect 22940 13462 22968 14486
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 22940 12714 22968 13398
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 22928 12708 22980 12714
rect 22928 12650 22980 12656
rect 22940 12102 22968 12650
rect 22928 12096 22980 12102
rect 22928 12038 22980 12044
rect 22940 11694 22968 12038
rect 23032 11801 23060 12718
rect 23018 11792 23074 11801
rect 23018 11727 23074 11736
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22836 9988 22888 9994
rect 22836 9930 22888 9936
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22560 9172 22612 9178
rect 22560 9114 22612 9120
rect 22572 8634 22600 9114
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22664 8362 22692 9318
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22756 8566 22784 8978
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22926 8528 22982 8537
rect 22926 8463 22982 8472
rect 22940 8430 22968 8463
rect 22928 8424 22980 8430
rect 22928 8366 22980 8372
rect 22192 8356 22244 8362
rect 22192 8298 22244 8304
rect 22652 8356 22704 8362
rect 22652 8298 22704 8304
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 21640 8016 21692 8022
rect 21640 7958 21692 7964
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21928 7342 21956 8026
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 21916 7336 21968 7342
rect 21916 7278 21968 7284
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 22940 4282 22968 8366
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 23032 3913 23060 4014
rect 23018 3904 23074 3913
rect 4322 3836 4630 3845
rect 23018 3839 23074 3848
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
<< via2 >>
rect 4328 23418 4384 23420
rect 4408 23418 4464 23420
rect 4488 23418 4544 23420
rect 4568 23418 4624 23420
rect 4328 23366 4374 23418
rect 4374 23366 4384 23418
rect 4408 23366 4438 23418
rect 4438 23366 4450 23418
rect 4450 23366 4464 23418
rect 4488 23366 4502 23418
rect 4502 23366 4514 23418
rect 4514 23366 4544 23418
rect 4568 23366 4578 23418
rect 4578 23366 4624 23418
rect 4328 23364 4384 23366
rect 4408 23364 4464 23366
rect 4488 23364 4544 23366
rect 4568 23364 4624 23366
rect 3668 22874 3724 22876
rect 3748 22874 3804 22876
rect 3828 22874 3884 22876
rect 3908 22874 3964 22876
rect 3668 22822 3714 22874
rect 3714 22822 3724 22874
rect 3748 22822 3778 22874
rect 3778 22822 3790 22874
rect 3790 22822 3804 22874
rect 3828 22822 3842 22874
rect 3842 22822 3854 22874
rect 3854 22822 3884 22874
rect 3908 22822 3918 22874
rect 3918 22822 3964 22874
rect 3668 22820 3724 22822
rect 3748 22820 3804 22822
rect 3828 22820 3884 22822
rect 3908 22820 3964 22822
rect 4328 22330 4384 22332
rect 4408 22330 4464 22332
rect 4488 22330 4544 22332
rect 4568 22330 4624 22332
rect 4328 22278 4374 22330
rect 4374 22278 4384 22330
rect 4408 22278 4438 22330
rect 4438 22278 4450 22330
rect 4450 22278 4464 22330
rect 4488 22278 4502 22330
rect 4502 22278 4514 22330
rect 4514 22278 4544 22330
rect 4568 22278 4578 22330
rect 4578 22278 4624 22330
rect 4328 22276 4384 22278
rect 4408 22276 4464 22278
rect 4488 22276 4544 22278
rect 4568 22276 4624 22278
rect 3668 21786 3724 21788
rect 3748 21786 3804 21788
rect 3828 21786 3884 21788
rect 3908 21786 3964 21788
rect 3668 21734 3714 21786
rect 3714 21734 3724 21786
rect 3748 21734 3778 21786
rect 3778 21734 3790 21786
rect 3790 21734 3804 21786
rect 3828 21734 3842 21786
rect 3842 21734 3854 21786
rect 3854 21734 3884 21786
rect 3908 21734 3918 21786
rect 3918 21734 3964 21786
rect 3668 21732 3724 21734
rect 3748 21732 3804 21734
rect 3828 21732 3884 21734
rect 3908 21732 3964 21734
rect 4328 21242 4384 21244
rect 4408 21242 4464 21244
rect 4488 21242 4544 21244
rect 4568 21242 4624 21244
rect 4328 21190 4374 21242
rect 4374 21190 4384 21242
rect 4408 21190 4438 21242
rect 4438 21190 4450 21242
rect 4450 21190 4464 21242
rect 4488 21190 4502 21242
rect 4502 21190 4514 21242
rect 4514 21190 4544 21242
rect 4568 21190 4578 21242
rect 4578 21190 4624 21242
rect 4328 21188 4384 21190
rect 4408 21188 4464 21190
rect 4488 21188 4544 21190
rect 4568 21188 4624 21190
rect 3668 20698 3724 20700
rect 3748 20698 3804 20700
rect 3828 20698 3884 20700
rect 3908 20698 3964 20700
rect 3668 20646 3714 20698
rect 3714 20646 3724 20698
rect 3748 20646 3778 20698
rect 3778 20646 3790 20698
rect 3790 20646 3804 20698
rect 3828 20646 3842 20698
rect 3842 20646 3854 20698
rect 3854 20646 3884 20698
rect 3908 20646 3918 20698
rect 3918 20646 3964 20698
rect 3668 20644 3724 20646
rect 3748 20644 3804 20646
rect 3828 20644 3884 20646
rect 3908 20644 3964 20646
rect 4328 20154 4384 20156
rect 4408 20154 4464 20156
rect 4488 20154 4544 20156
rect 4568 20154 4624 20156
rect 4328 20102 4374 20154
rect 4374 20102 4384 20154
rect 4408 20102 4438 20154
rect 4438 20102 4450 20154
rect 4450 20102 4464 20154
rect 4488 20102 4502 20154
rect 4502 20102 4514 20154
rect 4514 20102 4544 20154
rect 4568 20102 4578 20154
rect 4578 20102 4624 20154
rect 4328 20100 4384 20102
rect 4408 20100 4464 20102
rect 4488 20100 4544 20102
rect 4568 20100 4624 20102
rect 3668 19610 3724 19612
rect 3748 19610 3804 19612
rect 3828 19610 3884 19612
rect 3908 19610 3964 19612
rect 3668 19558 3714 19610
rect 3714 19558 3724 19610
rect 3748 19558 3778 19610
rect 3778 19558 3790 19610
rect 3790 19558 3804 19610
rect 3828 19558 3842 19610
rect 3842 19558 3854 19610
rect 3854 19558 3884 19610
rect 3908 19558 3918 19610
rect 3918 19558 3964 19610
rect 3668 19556 3724 19558
rect 3748 19556 3804 19558
rect 3828 19556 3884 19558
rect 3908 19556 3964 19558
rect 4328 19066 4384 19068
rect 4408 19066 4464 19068
rect 4488 19066 4544 19068
rect 4568 19066 4624 19068
rect 4328 19014 4374 19066
rect 4374 19014 4384 19066
rect 4408 19014 4438 19066
rect 4438 19014 4450 19066
rect 4450 19014 4464 19066
rect 4488 19014 4502 19066
rect 4502 19014 4514 19066
rect 4514 19014 4544 19066
rect 4568 19014 4578 19066
rect 4578 19014 4624 19066
rect 4328 19012 4384 19014
rect 4408 19012 4464 19014
rect 4488 19012 4544 19014
rect 4568 19012 4624 19014
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 4328 17978 4384 17980
rect 4408 17978 4464 17980
rect 4488 17978 4544 17980
rect 4568 17978 4624 17980
rect 4328 17926 4374 17978
rect 4374 17926 4384 17978
rect 4408 17926 4438 17978
rect 4438 17926 4450 17978
rect 4450 17926 4464 17978
rect 4488 17926 4502 17978
rect 4502 17926 4514 17978
rect 4514 17926 4544 17978
rect 4568 17926 4578 17978
rect 4578 17926 4624 17978
rect 4328 17924 4384 17926
rect 4408 17924 4464 17926
rect 4488 17924 4544 17926
rect 4568 17924 4624 17926
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 4328 16890 4384 16892
rect 4408 16890 4464 16892
rect 4488 16890 4544 16892
rect 4568 16890 4624 16892
rect 4328 16838 4374 16890
rect 4374 16838 4384 16890
rect 4408 16838 4438 16890
rect 4438 16838 4450 16890
rect 4450 16838 4464 16890
rect 4488 16838 4502 16890
rect 4502 16838 4514 16890
rect 4514 16838 4544 16890
rect 4568 16838 4578 16890
rect 4578 16838 4624 16890
rect 4328 16836 4384 16838
rect 4408 16836 4464 16838
rect 4488 16836 4544 16838
rect 4568 16836 4624 16838
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 4328 15802 4384 15804
rect 4408 15802 4464 15804
rect 4488 15802 4544 15804
rect 4568 15802 4624 15804
rect 4328 15750 4374 15802
rect 4374 15750 4384 15802
rect 4408 15750 4438 15802
rect 4438 15750 4450 15802
rect 4450 15750 4464 15802
rect 4488 15750 4502 15802
rect 4502 15750 4514 15802
rect 4514 15750 4544 15802
rect 4568 15750 4578 15802
rect 4578 15750 4624 15802
rect 4328 15748 4384 15750
rect 4408 15748 4464 15750
rect 4488 15748 4544 15750
rect 4568 15748 4624 15750
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 4328 14714 4384 14716
rect 4408 14714 4464 14716
rect 4488 14714 4544 14716
rect 4568 14714 4624 14716
rect 4328 14662 4374 14714
rect 4374 14662 4384 14714
rect 4408 14662 4438 14714
rect 4438 14662 4450 14714
rect 4450 14662 4464 14714
rect 4488 14662 4502 14714
rect 4502 14662 4514 14714
rect 4514 14662 4544 14714
rect 4568 14662 4578 14714
rect 4578 14662 4624 14714
rect 4328 14660 4384 14662
rect 4408 14660 4464 14662
rect 4488 14660 4544 14662
rect 4568 14660 4624 14662
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 4328 13626 4384 13628
rect 4408 13626 4464 13628
rect 4488 13626 4544 13628
rect 4568 13626 4624 13628
rect 4328 13574 4374 13626
rect 4374 13574 4384 13626
rect 4408 13574 4438 13626
rect 4438 13574 4450 13626
rect 4450 13574 4464 13626
rect 4488 13574 4502 13626
rect 4502 13574 4514 13626
rect 4514 13574 4544 13626
rect 4568 13574 4578 13626
rect 4578 13574 4624 13626
rect 4328 13572 4384 13574
rect 4408 13572 4464 13574
rect 4488 13572 4544 13574
rect 4568 13572 4624 13574
rect 6642 18708 6644 18728
rect 6644 18708 6696 18728
rect 6696 18708 6698 18728
rect 6642 18672 6698 18708
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 4328 12538 4384 12540
rect 4408 12538 4464 12540
rect 4488 12538 4544 12540
rect 4568 12538 4624 12540
rect 4328 12486 4374 12538
rect 4374 12486 4384 12538
rect 4408 12486 4438 12538
rect 4438 12486 4450 12538
rect 4450 12486 4464 12538
rect 4488 12486 4502 12538
rect 4502 12486 4514 12538
rect 4514 12486 4544 12538
rect 4568 12486 4578 12538
rect 4578 12486 4624 12538
rect 4328 12484 4384 12486
rect 4408 12484 4464 12486
rect 4488 12484 4544 12486
rect 4568 12484 4624 12486
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 4328 11450 4384 11452
rect 4408 11450 4464 11452
rect 4488 11450 4544 11452
rect 4568 11450 4624 11452
rect 4328 11398 4374 11450
rect 4374 11398 4384 11450
rect 4408 11398 4438 11450
rect 4438 11398 4450 11450
rect 4450 11398 4464 11450
rect 4488 11398 4502 11450
rect 4502 11398 4514 11450
rect 4514 11398 4544 11450
rect 4568 11398 4578 11450
rect 4578 11398 4624 11450
rect 4328 11396 4384 11398
rect 4408 11396 4464 11398
rect 4488 11396 4544 11398
rect 4568 11396 4624 11398
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 4328 10362 4384 10364
rect 4408 10362 4464 10364
rect 4488 10362 4544 10364
rect 4568 10362 4624 10364
rect 4328 10310 4374 10362
rect 4374 10310 4384 10362
rect 4408 10310 4438 10362
rect 4438 10310 4450 10362
rect 4450 10310 4464 10362
rect 4488 10310 4502 10362
rect 4502 10310 4514 10362
rect 4514 10310 4544 10362
rect 4568 10310 4578 10362
rect 4578 10310 4624 10362
rect 4328 10308 4384 10310
rect 4408 10308 4464 10310
rect 4488 10308 4544 10310
rect 4568 10308 4624 10310
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 12070 21936 12126 21992
rect 12070 18844 12072 18864
rect 12072 18844 12124 18864
rect 12124 18844 12126 18864
rect 12070 18808 12126 18844
rect 14094 21936 14150 21992
rect 14186 20712 14242 20768
rect 14738 21428 14740 21448
rect 14740 21428 14792 21448
rect 14792 21428 14794 21448
rect 14738 21392 14794 21428
rect 15382 22344 15438 22400
rect 15014 18400 15070 18456
rect 14922 16516 14978 16552
rect 14922 16496 14924 16516
rect 14924 16496 14976 16516
rect 14976 16496 14978 16516
rect 16486 22344 16542 22400
rect 16578 21392 16634 21448
rect 18878 21428 18880 21448
rect 18880 21428 18932 21448
rect 18932 21428 18934 21448
rect 18878 21392 18934 21428
rect 16394 18844 16396 18864
rect 16396 18844 16448 18864
rect 16448 18844 16450 18864
rect 16394 18808 16450 18844
rect 15474 18672 15530 18728
rect 16394 18400 16450 18456
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 20074 8472 20130 8528
rect 19890 8336 19946 8392
rect 23018 19624 23074 19680
rect 21822 8336 21878 8392
rect 23018 11736 23074 11792
rect 22926 8472 22982 8528
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 23018 3848 23074 3904
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
<< metal3 >>
rect 4318 23424 4634 23425
rect 4318 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4634 23424
rect 4318 23359 4634 23360
rect 3658 22880 3974 22881
rect 3658 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3974 22880
rect 3658 22815 3974 22816
rect 15377 22402 15443 22405
rect 16481 22402 16547 22405
rect 15377 22400 16547 22402
rect 15377 22344 15382 22400
rect 15438 22344 16486 22400
rect 16542 22344 16547 22400
rect 15377 22342 16547 22344
rect 15377 22339 15443 22342
rect 16481 22339 16547 22342
rect 4318 22336 4634 22337
rect 4318 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4634 22336
rect 4318 22271 4634 22272
rect 12065 21994 12131 21997
rect 14089 21994 14155 21997
rect 12065 21992 14155 21994
rect 12065 21936 12070 21992
rect 12126 21936 14094 21992
rect 14150 21936 14155 21992
rect 12065 21934 14155 21936
rect 12065 21931 12131 21934
rect 14089 21931 14155 21934
rect 3658 21792 3974 21793
rect 3658 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3974 21792
rect 3658 21727 3974 21728
rect 14733 21450 14799 21453
rect 16573 21450 16639 21453
rect 18873 21450 18939 21453
rect 14733 21448 18939 21450
rect 14733 21392 14738 21448
rect 14794 21392 16578 21448
rect 16634 21392 18878 21448
rect 18934 21392 18939 21448
rect 14733 21390 18939 21392
rect 14733 21387 14799 21390
rect 16573 21387 16639 21390
rect 18873 21387 18939 21390
rect 4318 21248 4634 21249
rect 4318 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4634 21248
rect 4318 21183 4634 21184
rect 14181 20770 14247 20773
rect 14774 20770 14780 20772
rect 14181 20768 14780 20770
rect 14181 20712 14186 20768
rect 14242 20712 14780 20768
rect 14181 20710 14780 20712
rect 14181 20707 14247 20710
rect 14774 20708 14780 20710
rect 14844 20708 14850 20772
rect 3658 20704 3974 20705
rect 3658 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3974 20704
rect 3658 20639 3974 20640
rect 4318 20160 4634 20161
rect 4318 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4634 20160
rect 4318 20095 4634 20096
rect 23013 19682 23079 19685
rect 23600 19682 24000 19712
rect 23013 19680 24000 19682
rect 23013 19624 23018 19680
rect 23074 19624 24000 19680
rect 23013 19622 24000 19624
rect 23013 19619 23079 19622
rect 3658 19616 3974 19617
rect 3658 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3974 19616
rect 23600 19592 24000 19622
rect 3658 19551 3974 19552
rect 4318 19072 4634 19073
rect 4318 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4634 19072
rect 4318 19007 4634 19008
rect 12065 18866 12131 18869
rect 16389 18866 16455 18869
rect 12065 18864 16455 18866
rect 12065 18808 12070 18864
rect 12126 18808 16394 18864
rect 16450 18808 16455 18864
rect 12065 18806 16455 18808
rect 12065 18803 12131 18806
rect 16389 18803 16455 18806
rect 6637 18730 6703 18733
rect 15469 18730 15535 18733
rect 6637 18728 15535 18730
rect 6637 18672 6642 18728
rect 6698 18672 15474 18728
rect 15530 18672 15535 18728
rect 6637 18670 15535 18672
rect 6637 18667 6703 18670
rect 15469 18667 15535 18670
rect 3658 18528 3974 18529
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 15009 18458 15075 18461
rect 16389 18458 16455 18461
rect 15009 18456 16455 18458
rect 15009 18400 15014 18456
rect 15070 18400 16394 18456
rect 16450 18400 16455 18456
rect 15009 18398 16455 18400
rect 15009 18395 15075 18398
rect 16389 18395 16455 18398
rect 4318 17984 4634 17985
rect 4318 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4634 17984
rect 4318 17919 4634 17920
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 4318 16896 4634 16897
rect 4318 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4634 16896
rect 4318 16831 4634 16832
rect 14774 16492 14780 16556
rect 14844 16554 14850 16556
rect 14917 16554 14983 16557
rect 14844 16552 14983 16554
rect 14844 16496 14922 16552
rect 14978 16496 14983 16552
rect 14844 16494 14983 16496
rect 14844 16492 14850 16494
rect 14917 16491 14983 16494
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 4318 15808 4634 15809
rect 4318 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4634 15808
rect 4318 15743 4634 15744
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 4318 14720 4634 14721
rect 4318 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4634 14720
rect 4318 14655 4634 14656
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 4318 13632 4634 13633
rect 4318 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4634 13632
rect 4318 13567 4634 13568
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 4318 12544 4634 12545
rect 4318 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4634 12544
rect 4318 12479 4634 12480
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 23013 11794 23079 11797
rect 23600 11794 24000 11824
rect 23013 11792 24000 11794
rect 23013 11736 23018 11792
rect 23074 11736 24000 11792
rect 23013 11734 24000 11736
rect 23013 11731 23079 11734
rect 23600 11704 24000 11734
rect 4318 11456 4634 11457
rect 4318 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4634 11456
rect 4318 11391 4634 11392
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 4318 10368 4634 10369
rect 4318 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4634 10368
rect 4318 10303 4634 10304
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 20069 8530 20135 8533
rect 22921 8530 22987 8533
rect 20069 8528 22987 8530
rect 20069 8472 20074 8528
rect 20130 8472 22926 8528
rect 22982 8472 22987 8528
rect 20069 8470 22987 8472
rect 20069 8467 20135 8470
rect 22921 8467 22987 8470
rect 19885 8394 19951 8397
rect 21817 8394 21883 8397
rect 19885 8392 21883 8394
rect 19885 8336 19890 8392
rect 19946 8336 21822 8392
rect 21878 8336 21883 8392
rect 19885 8334 21883 8336
rect 19885 8331 19951 8334
rect 21817 8331 21883 8334
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 23013 3906 23079 3909
rect 23600 3906 24000 3936
rect 23013 3904 24000 3906
rect 23013 3848 23018 3904
rect 23074 3848 24000 3904
rect 23013 3846 24000 3848
rect 23013 3843 23079 3846
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 23600 3816 24000 3846
rect 4318 3775 4634 3776
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
<< via3 >>
rect 4324 23420 4388 23424
rect 4324 23364 4328 23420
rect 4328 23364 4384 23420
rect 4384 23364 4388 23420
rect 4324 23360 4388 23364
rect 4404 23420 4468 23424
rect 4404 23364 4408 23420
rect 4408 23364 4464 23420
rect 4464 23364 4468 23420
rect 4404 23360 4468 23364
rect 4484 23420 4548 23424
rect 4484 23364 4488 23420
rect 4488 23364 4544 23420
rect 4544 23364 4548 23420
rect 4484 23360 4548 23364
rect 4564 23420 4628 23424
rect 4564 23364 4568 23420
rect 4568 23364 4624 23420
rect 4624 23364 4628 23420
rect 4564 23360 4628 23364
rect 3664 22876 3728 22880
rect 3664 22820 3668 22876
rect 3668 22820 3724 22876
rect 3724 22820 3728 22876
rect 3664 22816 3728 22820
rect 3744 22876 3808 22880
rect 3744 22820 3748 22876
rect 3748 22820 3804 22876
rect 3804 22820 3808 22876
rect 3744 22816 3808 22820
rect 3824 22876 3888 22880
rect 3824 22820 3828 22876
rect 3828 22820 3884 22876
rect 3884 22820 3888 22876
rect 3824 22816 3888 22820
rect 3904 22876 3968 22880
rect 3904 22820 3908 22876
rect 3908 22820 3964 22876
rect 3964 22820 3968 22876
rect 3904 22816 3968 22820
rect 4324 22332 4388 22336
rect 4324 22276 4328 22332
rect 4328 22276 4384 22332
rect 4384 22276 4388 22332
rect 4324 22272 4388 22276
rect 4404 22332 4468 22336
rect 4404 22276 4408 22332
rect 4408 22276 4464 22332
rect 4464 22276 4468 22332
rect 4404 22272 4468 22276
rect 4484 22332 4548 22336
rect 4484 22276 4488 22332
rect 4488 22276 4544 22332
rect 4544 22276 4548 22332
rect 4484 22272 4548 22276
rect 4564 22332 4628 22336
rect 4564 22276 4568 22332
rect 4568 22276 4624 22332
rect 4624 22276 4628 22332
rect 4564 22272 4628 22276
rect 3664 21788 3728 21792
rect 3664 21732 3668 21788
rect 3668 21732 3724 21788
rect 3724 21732 3728 21788
rect 3664 21728 3728 21732
rect 3744 21788 3808 21792
rect 3744 21732 3748 21788
rect 3748 21732 3804 21788
rect 3804 21732 3808 21788
rect 3744 21728 3808 21732
rect 3824 21788 3888 21792
rect 3824 21732 3828 21788
rect 3828 21732 3884 21788
rect 3884 21732 3888 21788
rect 3824 21728 3888 21732
rect 3904 21788 3968 21792
rect 3904 21732 3908 21788
rect 3908 21732 3964 21788
rect 3964 21732 3968 21788
rect 3904 21728 3968 21732
rect 4324 21244 4388 21248
rect 4324 21188 4328 21244
rect 4328 21188 4384 21244
rect 4384 21188 4388 21244
rect 4324 21184 4388 21188
rect 4404 21244 4468 21248
rect 4404 21188 4408 21244
rect 4408 21188 4464 21244
rect 4464 21188 4468 21244
rect 4404 21184 4468 21188
rect 4484 21244 4548 21248
rect 4484 21188 4488 21244
rect 4488 21188 4544 21244
rect 4544 21188 4548 21244
rect 4484 21184 4548 21188
rect 4564 21244 4628 21248
rect 4564 21188 4568 21244
rect 4568 21188 4624 21244
rect 4624 21188 4628 21244
rect 4564 21184 4628 21188
rect 14780 20708 14844 20772
rect 3664 20700 3728 20704
rect 3664 20644 3668 20700
rect 3668 20644 3724 20700
rect 3724 20644 3728 20700
rect 3664 20640 3728 20644
rect 3744 20700 3808 20704
rect 3744 20644 3748 20700
rect 3748 20644 3804 20700
rect 3804 20644 3808 20700
rect 3744 20640 3808 20644
rect 3824 20700 3888 20704
rect 3824 20644 3828 20700
rect 3828 20644 3884 20700
rect 3884 20644 3888 20700
rect 3824 20640 3888 20644
rect 3904 20700 3968 20704
rect 3904 20644 3908 20700
rect 3908 20644 3964 20700
rect 3964 20644 3968 20700
rect 3904 20640 3968 20644
rect 4324 20156 4388 20160
rect 4324 20100 4328 20156
rect 4328 20100 4384 20156
rect 4384 20100 4388 20156
rect 4324 20096 4388 20100
rect 4404 20156 4468 20160
rect 4404 20100 4408 20156
rect 4408 20100 4464 20156
rect 4464 20100 4468 20156
rect 4404 20096 4468 20100
rect 4484 20156 4548 20160
rect 4484 20100 4488 20156
rect 4488 20100 4544 20156
rect 4544 20100 4548 20156
rect 4484 20096 4548 20100
rect 4564 20156 4628 20160
rect 4564 20100 4568 20156
rect 4568 20100 4624 20156
rect 4624 20100 4628 20156
rect 4564 20096 4628 20100
rect 3664 19612 3728 19616
rect 3664 19556 3668 19612
rect 3668 19556 3724 19612
rect 3724 19556 3728 19612
rect 3664 19552 3728 19556
rect 3744 19612 3808 19616
rect 3744 19556 3748 19612
rect 3748 19556 3804 19612
rect 3804 19556 3808 19612
rect 3744 19552 3808 19556
rect 3824 19612 3888 19616
rect 3824 19556 3828 19612
rect 3828 19556 3884 19612
rect 3884 19556 3888 19612
rect 3824 19552 3888 19556
rect 3904 19612 3968 19616
rect 3904 19556 3908 19612
rect 3908 19556 3964 19612
rect 3964 19556 3968 19612
rect 3904 19552 3968 19556
rect 4324 19068 4388 19072
rect 4324 19012 4328 19068
rect 4328 19012 4384 19068
rect 4384 19012 4388 19068
rect 4324 19008 4388 19012
rect 4404 19068 4468 19072
rect 4404 19012 4408 19068
rect 4408 19012 4464 19068
rect 4464 19012 4468 19068
rect 4404 19008 4468 19012
rect 4484 19068 4548 19072
rect 4484 19012 4488 19068
rect 4488 19012 4544 19068
rect 4544 19012 4548 19068
rect 4484 19008 4548 19012
rect 4564 19068 4628 19072
rect 4564 19012 4568 19068
rect 4568 19012 4624 19068
rect 4624 19012 4628 19068
rect 4564 19008 4628 19012
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 4324 17980 4388 17984
rect 4324 17924 4328 17980
rect 4328 17924 4384 17980
rect 4384 17924 4388 17980
rect 4324 17920 4388 17924
rect 4404 17980 4468 17984
rect 4404 17924 4408 17980
rect 4408 17924 4464 17980
rect 4464 17924 4468 17980
rect 4404 17920 4468 17924
rect 4484 17980 4548 17984
rect 4484 17924 4488 17980
rect 4488 17924 4544 17980
rect 4544 17924 4548 17980
rect 4484 17920 4548 17924
rect 4564 17980 4628 17984
rect 4564 17924 4568 17980
rect 4568 17924 4624 17980
rect 4624 17924 4628 17980
rect 4564 17920 4628 17924
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 4324 16892 4388 16896
rect 4324 16836 4328 16892
rect 4328 16836 4384 16892
rect 4384 16836 4388 16892
rect 4324 16832 4388 16836
rect 4404 16892 4468 16896
rect 4404 16836 4408 16892
rect 4408 16836 4464 16892
rect 4464 16836 4468 16892
rect 4404 16832 4468 16836
rect 4484 16892 4548 16896
rect 4484 16836 4488 16892
rect 4488 16836 4544 16892
rect 4544 16836 4548 16892
rect 4484 16832 4548 16836
rect 4564 16892 4628 16896
rect 4564 16836 4568 16892
rect 4568 16836 4624 16892
rect 4624 16836 4628 16892
rect 4564 16832 4628 16836
rect 14780 16492 14844 16556
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 4324 15804 4388 15808
rect 4324 15748 4328 15804
rect 4328 15748 4384 15804
rect 4384 15748 4388 15804
rect 4324 15744 4388 15748
rect 4404 15804 4468 15808
rect 4404 15748 4408 15804
rect 4408 15748 4464 15804
rect 4464 15748 4468 15804
rect 4404 15744 4468 15748
rect 4484 15804 4548 15808
rect 4484 15748 4488 15804
rect 4488 15748 4544 15804
rect 4544 15748 4548 15804
rect 4484 15744 4548 15748
rect 4564 15804 4628 15808
rect 4564 15748 4568 15804
rect 4568 15748 4624 15804
rect 4624 15748 4628 15804
rect 4564 15744 4628 15748
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 4324 14716 4388 14720
rect 4324 14660 4328 14716
rect 4328 14660 4384 14716
rect 4384 14660 4388 14716
rect 4324 14656 4388 14660
rect 4404 14716 4468 14720
rect 4404 14660 4408 14716
rect 4408 14660 4464 14716
rect 4464 14660 4468 14716
rect 4404 14656 4468 14660
rect 4484 14716 4548 14720
rect 4484 14660 4488 14716
rect 4488 14660 4544 14716
rect 4544 14660 4548 14716
rect 4484 14656 4548 14660
rect 4564 14716 4628 14720
rect 4564 14660 4568 14716
rect 4568 14660 4624 14716
rect 4624 14660 4628 14716
rect 4564 14656 4628 14660
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 4324 13628 4388 13632
rect 4324 13572 4328 13628
rect 4328 13572 4384 13628
rect 4384 13572 4388 13628
rect 4324 13568 4388 13572
rect 4404 13628 4468 13632
rect 4404 13572 4408 13628
rect 4408 13572 4464 13628
rect 4464 13572 4468 13628
rect 4404 13568 4468 13572
rect 4484 13628 4548 13632
rect 4484 13572 4488 13628
rect 4488 13572 4544 13628
rect 4544 13572 4548 13628
rect 4484 13568 4548 13572
rect 4564 13628 4628 13632
rect 4564 13572 4568 13628
rect 4568 13572 4624 13628
rect 4624 13572 4628 13628
rect 4564 13568 4628 13572
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 4324 12540 4388 12544
rect 4324 12484 4328 12540
rect 4328 12484 4384 12540
rect 4384 12484 4388 12540
rect 4324 12480 4388 12484
rect 4404 12540 4468 12544
rect 4404 12484 4408 12540
rect 4408 12484 4464 12540
rect 4464 12484 4468 12540
rect 4404 12480 4468 12484
rect 4484 12540 4548 12544
rect 4484 12484 4488 12540
rect 4488 12484 4544 12540
rect 4544 12484 4548 12540
rect 4484 12480 4548 12484
rect 4564 12540 4628 12544
rect 4564 12484 4568 12540
rect 4568 12484 4624 12540
rect 4624 12484 4628 12540
rect 4564 12480 4628 12484
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 4324 11452 4388 11456
rect 4324 11396 4328 11452
rect 4328 11396 4384 11452
rect 4384 11396 4388 11452
rect 4324 11392 4388 11396
rect 4404 11452 4468 11456
rect 4404 11396 4408 11452
rect 4408 11396 4464 11452
rect 4464 11396 4468 11452
rect 4404 11392 4468 11396
rect 4484 11452 4548 11456
rect 4484 11396 4488 11452
rect 4488 11396 4544 11452
rect 4544 11396 4548 11452
rect 4484 11392 4548 11396
rect 4564 11452 4628 11456
rect 4564 11396 4568 11452
rect 4568 11396 4624 11452
rect 4624 11396 4628 11452
rect 4564 11392 4628 11396
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 4324 10364 4388 10368
rect 4324 10308 4328 10364
rect 4328 10308 4384 10364
rect 4384 10308 4388 10364
rect 4324 10304 4388 10308
rect 4404 10364 4468 10368
rect 4404 10308 4408 10364
rect 4408 10308 4464 10364
rect 4464 10308 4468 10364
rect 4404 10304 4468 10308
rect 4484 10364 4548 10368
rect 4484 10308 4488 10364
rect 4488 10308 4544 10364
rect 4544 10308 4548 10364
rect 4484 10304 4548 10308
rect 4564 10364 4628 10368
rect 4564 10308 4568 10364
rect 4568 10308 4624 10364
rect 4624 10308 4628 10364
rect 4564 10304 4628 10308
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
<< metal4 >>
rect 3656 22880 3976 23440
rect 3656 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3976 22880
rect 3656 21792 3976 22816
rect 3656 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3976 21792
rect 3656 20704 3976 21728
rect 3656 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3976 20704
rect 3656 19616 3976 20640
rect 3656 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3976 19616
rect 3656 18528 3976 19552
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 3656 17440 3976 18464
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3656 15264 3976 16288
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3656 14176 3976 15200
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3656 12000 3976 13024
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 23424 4636 23440
rect 4316 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4636 23424
rect 4316 22336 4636 23360
rect 4316 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4636 22336
rect 4316 21248 4636 22272
rect 4316 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4636 21248
rect 4316 20160 4636 21184
rect 14779 20772 14845 20773
rect 14779 20708 14780 20772
rect 14844 20708 14845 20772
rect 14779 20707 14845 20708
rect 4316 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4636 20160
rect 4316 19072 4636 20096
rect 4316 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4636 19072
rect 4316 17984 4636 19008
rect 4316 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4636 17984
rect 4316 16896 4636 17920
rect 4316 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4636 16896
rect 4316 15808 4636 16832
rect 14782 16557 14842 20707
rect 14779 16556 14845 16557
rect 14779 16492 14780 16556
rect 14844 16492 14845 16556
rect 14779 16491 14845 16492
rect 4316 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4636 15808
rect 4316 14720 4636 15744
rect 4316 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4636 14720
rect 4316 13632 4636 14656
rect 4316 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4636 13632
rect 4316 12544 4636 13568
rect 4316 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4636 12544
rect 4316 11456 4636 12480
rect 4316 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4636 11456
rect 4316 10368 4636 11392
rect 4316 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4636 10368
rect 4316 9280 4636 10304
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
use sky130_fd_sc_hd__inv_2  _0490_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 23000 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1723858470
transform 1 0 20976 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1723858470
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1723858470
transform -1 0 4600 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1723858470
transform 1 0 8372 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_6  _0495_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 20424 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0496_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6348 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0497_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6440 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0498_
timestamp 1723858470
transform 1 0 8924 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0499_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10212 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0500_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0501_
timestamp 1723858470
transform 1 0 12512 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0502_
timestamp 1723858470
transform 1 0 14260 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0503_
timestamp 1723858470
transform 1 0 16100 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0504_
timestamp 1723858470
transform 1 0 16928 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0505_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 17940 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0506_
timestamp 1723858470
transform 1 0 19320 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0507_
timestamp 1723858470
transform -1 0 20792 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0508_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21620 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0509_
timestamp 1723858470
transform 1 0 22172 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _0510_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0511_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5796 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0512_
timestamp 1723858470
transform 1 0 4692 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0513_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5244 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0514_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5060 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0515_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _0516_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4968 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0517_
timestamp 1723858470
transform 1 0 4968 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0518_
timestamp 1723858470
transform -1 0 5336 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0519_
timestamp 1723858470
transform 1 0 5796 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0520_
timestamp 1723858470
transform 1 0 4600 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0521_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5428 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0522_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5704 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0523_
timestamp 1723858470
transform 1 0 7176 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0524_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9476 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0525_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8832 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0526_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6256 0 1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__mux2_1  _0527_
timestamp 1723858470
transform 1 0 8372 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0528_
timestamp 1723858470
transform 1 0 7452 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _0529_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4876 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0530_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5888 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0531_
timestamp 1723858470
transform 1 0 7544 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0532_
timestamp 1723858470
transform 1 0 10120 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0533_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9292 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0534_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9660 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0535_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 10764 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0536_
timestamp 1723858470
transform -1 0 9016 0 -1 21216
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0537_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8832 0 -1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_2  _0538_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4600 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _0539_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6532 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0540_
timestamp 1723858470
transform 1 0 8372 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0541_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7176 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0542_
timestamp 1723858470
transform 1 0 9568 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0543_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8188 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0544_
timestamp 1723858470
transform 1 0 9844 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0545_
timestamp 1723858470
transform -1 0 9844 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0546_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9292 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0547_
timestamp 1723858470
transform 1 0 8648 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0548_
timestamp 1723858470
transform 1 0 8648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0549_
timestamp 1723858470
transform -1 0 9476 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1723858470
transform 1 0 10212 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0551_
timestamp 1723858470
transform 1 0 8924 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0552_
timestamp 1723858470
transform -1 0 9660 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0553_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 10396 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0554_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 12052 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0555_
timestamp 1723858470
transform -1 0 12972 0 1 19040
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1723858470
transform 1 0 10212 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0557_
timestamp 1723858470
transform 1 0 5980 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0558_
timestamp 1723858470
transform 1 0 5428 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_2  _0559_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6440 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0560_
timestamp 1723858470
transform -1 0 7084 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0561_
timestamp 1723858470
transform 1 0 6532 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0562_
timestamp 1723858470
transform -1 0 10580 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0563_
timestamp 1723858470
transform -1 0 9200 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0564_
timestamp 1723858470
transform 1 0 9844 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0565_
timestamp 1723858470
transform -1 0 9936 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0566_
timestamp 1723858470
transform -1 0 10028 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0567_
timestamp 1723858470
transform 1 0 10028 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0568_
timestamp 1723858470
transform 1 0 8740 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0569_
timestamp 1723858470
transform 1 0 9016 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0570_
timestamp 1723858470
transform 1 0 9384 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _0571_
timestamp 1723858470
transform -1 0 10948 0 1 19040
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0572_
timestamp 1723858470
transform -1 0 10856 0 -1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_1  _0573_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4876 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0574_
timestamp 1723858470
transform -1 0 7084 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0575_
timestamp 1723858470
transform 1 0 5428 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0576_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7912 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0577_
timestamp 1723858470
transform 1 0 7084 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0578_
timestamp 1723858470
transform 1 0 6256 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0579_
timestamp 1723858470
transform 1 0 8372 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0580_
timestamp 1723858470
transform 1 0 9200 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0581_
timestamp 1723858470
transform 1 0 9568 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0582_
timestamp 1723858470
transform 1 0 9292 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0583_
timestamp 1723858470
transform 1 0 10764 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0584_
timestamp 1723858470
transform -1 0 10764 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0585_
timestamp 1723858470
transform 1 0 10856 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0586_
timestamp 1723858470
transform 1 0 10212 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0587_
timestamp 1723858470
transform -1 0 10856 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0588_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 10212 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0589_
timestamp 1723858470
transform 1 0 10212 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0590_
timestamp 1723858470
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _0591_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10948 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0592_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7544 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__o31a_1  _0593_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6440 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0594_
timestamp 1723858470
transform 1 0 5336 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0595_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6164 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0596_
timestamp 1723858470
transform 1 0 6164 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0597_
timestamp 1723858470
transform 1 0 5796 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0598_
timestamp 1723858470
transform 1 0 7636 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0599_
timestamp 1723858470
transform -1 0 7820 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _0600_
timestamp 1723858470
transform 1 0 8556 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0601_
timestamp 1723858470
transform 1 0 7912 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0602_
timestamp 1723858470
transform 1 0 12052 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0603_
timestamp 1723858470
transform 1 0 11040 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0604_
timestamp 1723858470
transform 1 0 11960 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0605_
timestamp 1723858470
transform 1 0 11684 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0606_
timestamp 1723858470
transform -1 0 11960 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0607_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9936 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0608_
timestamp 1723858470
transform 1 0 9844 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0609_
timestamp 1723858470
transform 1 0 10764 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _0610_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10948 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0611_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12052 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0612_
timestamp 1723858470
transform 1 0 11500 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0613_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 11592 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0614_
timestamp 1723858470
transform -1 0 16560 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0615_
timestamp 1723858470
transform 1 0 15088 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0616_
timestamp 1723858470
transform 1 0 16928 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0617_
timestamp 1723858470
transform -1 0 16192 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0618_
timestamp 1723858470
transform 1 0 16284 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0619_
timestamp 1723858470
transform -1 0 16192 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _0620_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 11040 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0621_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10856 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0622_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12788 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0623_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12236 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0624_
timestamp 1723858470
transform -1 0 12604 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0625_
timestamp 1723858470
transform -1 0 13432 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0626_
timestamp 1723858470
transform 1 0 6900 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0627_
timestamp 1723858470
transform 1 0 12972 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0628_
timestamp 1723858470
transform 1 0 11684 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0629_
timestamp 1723858470
transform 1 0 12328 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0630_
timestamp 1723858470
transform -1 0 13064 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0631_
timestamp 1723858470
transform 1 0 12696 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0632_
timestamp 1723858470
transform -1 0 13340 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0633_
timestamp 1723858470
transform -1 0 13616 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0634_
timestamp 1723858470
transform 1 0 12788 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2ai_1  _0635_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 12328 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0636_
timestamp 1723858470
transform -1 0 15180 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_4  _0637_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 16100 0 -1 22304
box -38 -48 1418 592
use sky130_fd_sc_hd__a21oi_2  _0638_
timestamp 1723858470
transform 1 0 18768 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0639_
timestamp 1723858470
transform 1 0 18124 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0640_
timestamp 1723858470
transform 1 0 19964 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0641_
timestamp 1723858470
transform -1 0 20332 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _0642_
timestamp 1723858470
transform -1 0 11684 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _0643_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12052 0 -1 22304
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0644_
timestamp 1723858470
transform -1 0 14536 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0645_
timestamp 1723858470
transform -1 0 13432 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0646_
timestamp 1723858470
transform -1 0 12880 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0647_
timestamp 1723858470
transform 1 0 13708 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0648_
timestamp 1723858470
transform -1 0 13432 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0649_
timestamp 1723858470
transform 1 0 14260 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0650_
timestamp 1723858470
transform 1 0 14260 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _0651_
timestamp 1723858470
transform -1 0 13892 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0652_
timestamp 1723858470
transform 1 0 14904 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0653_
timestamp 1723858470
transform -1 0 14904 0 -1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0654_
timestamp 1723858470
transform -1 0 14352 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0655_
timestamp 1723858470
transform 1 0 13708 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0656_
timestamp 1723858470
transform 1 0 14076 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0657_
timestamp 1723858470
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _0658_
timestamp 1723858470
transform 1 0 19044 0 -1 22304
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_1  _0659_
timestamp 1723858470
transform 1 0 10304 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0660_
timestamp 1723858470
transform 1 0 10120 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 1723858470
transform 1 0 10580 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0662_
timestamp 1723858470
transform 1 0 7544 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0663_
timestamp 1723858470
transform 1 0 9200 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0664_
timestamp 1723858470
transform 1 0 9108 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0665_
timestamp 1723858470
transform 1 0 10948 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_1  _0666_
timestamp 1723858470
transform 1 0 13524 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0667_
timestamp 1723858470
transform 1 0 14536 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0668_
timestamp 1723858470
transform 1 0 13616 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0669_
timestamp 1723858470
transform -1 0 15640 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0670_
timestamp 1723858470
transform -1 0 15640 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0671_
timestamp 1723858470
transform 1 0 14996 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0672_
timestamp 1723858470
transform -1 0 14904 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0673_
timestamp 1723858470
transform -1 0 14812 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0674_
timestamp 1723858470
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0675_
timestamp 1723858470
transform 1 0 14536 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0676_
timestamp 1723858470
transform 1 0 13524 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0677_
timestamp 1723858470
transform -1 0 8924 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0678_
timestamp 1723858470
transform 1 0 8464 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0679_
timestamp 1723858470
transform 1 0 11132 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0680_
timestamp 1723858470
transform -1 0 10948 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0681_
timestamp 1723858470
transform 1 0 12604 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0682_
timestamp 1723858470
transform 1 0 12236 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0683_
timestamp 1723858470
transform 1 0 13524 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0684_
timestamp 1723858470
transform 1 0 12972 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0685_
timestamp 1723858470
transform -1 0 15548 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0686_
timestamp 1723858470
transform 1 0 14076 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0687_
timestamp 1723858470
transform 1 0 13984 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0688_
timestamp 1723858470
transform -1 0 14996 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0689_
timestamp 1723858470
transform 1 0 14444 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1723858470
transform 1 0 14628 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0691_
timestamp 1723858470
transform 1 0 14536 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1723858470
transform 1 0 15364 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0693_
timestamp 1723858470
transform 1 0 9752 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0694_
timestamp 1723858470
transform 1 0 8924 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0695_
timestamp 1723858470
transform 1 0 10396 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0696_
timestamp 1723858470
transform 1 0 10764 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0697_
timestamp 1723858470
transform 1 0 12144 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0698_
timestamp 1723858470
transform -1 0 14076 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0699_
timestamp 1723858470
transform 1 0 13616 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0700_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 13984 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 1723858470
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0702_
timestamp 1723858470
transform -1 0 15732 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0703_
timestamp 1723858470
transform 1 0 14536 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1723858470
transform 1 0 16100 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0705_
timestamp 1723858470
transform 1 0 5060 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0706_
timestamp 1723858470
transform 1 0 5060 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0707_
timestamp 1723858470
transform 1 0 7912 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0708_
timestamp 1723858470
transform 1 0 6624 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0709_
timestamp 1723858470
transform 1 0 8096 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _0710_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9292 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0711_
timestamp 1723858470
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0712_
timestamp 1723858470
transform 1 0 10580 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0713_
timestamp 1723858470
transform 1 0 12512 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _0714_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12052 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0715_
timestamp 1723858470
transform 1 0 13800 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1723858470
transform 1 0 17296 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0717_
timestamp 1723858470
transform 1 0 13156 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0718_
timestamp 1723858470
transform 1 0 15180 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0719_
timestamp 1723858470
transform -1 0 14628 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0720_
timestamp 1723858470
transform -1 0 14536 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0721_
timestamp 1723858470
transform 1 0 15640 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0722_
timestamp 1723858470
transform 1 0 16100 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0723_
timestamp 1723858470
transform 1 0 16100 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 1723858470
transform 1 0 6900 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0725_
timestamp 1723858470
transform 1 0 6440 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0726_
timestamp 1723858470
transform 1 0 6624 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0727_
timestamp 1723858470
transform -1 0 6256 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0728_
timestamp 1723858470
transform 1 0 6808 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0729_
timestamp 1723858470
transform 1 0 6440 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0730_
timestamp 1723858470
transform 1 0 7636 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0731_
timestamp 1723858470
transform 1 0 6624 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0732_
timestamp 1723858470
transform 1 0 15824 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0733_
timestamp 1723858470
transform 1 0 15180 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0734_
timestamp 1723858470
transform -1 0 16744 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0735_
timestamp 1723858470
transform 1 0 11684 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0736_
timestamp 1723858470
transform 1 0 15548 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0737_
timestamp 1723858470
transform -1 0 17020 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0738_
timestamp 1723858470
transform 1 0 16100 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1723858470
transform 1 0 17020 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0740_
timestamp 1723858470
transform -1 0 17020 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0741_
timestamp 1723858470
transform -1 0 17388 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0742_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 16744 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1723858470
transform 1 0 16284 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0744_
timestamp 1723858470
transform 1 0 15548 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0745_
timestamp 1723858470
transform -1 0 17756 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0746_
timestamp 1723858470
transform 1 0 17572 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0747_
timestamp 1723858470
transform -1 0 17480 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0748_
timestamp 1723858470
transform -1 0 17940 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0749_
timestamp 1723858470
transform 1 0 7360 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0750_
timestamp 1723858470
transform 1 0 17572 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0751_
timestamp 1723858470
transform -1 0 17572 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0752_
timestamp 1723858470
transform -1 0 17204 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0753_
timestamp 1723858470
transform 1 0 17204 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0754_
timestamp 1723858470
transform -1 0 16652 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0755_
timestamp 1723858470
transform -1 0 18584 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0756_
timestamp 1723858470
transform 1 0 17848 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0757_
timestamp 1723858470
transform 1 0 18768 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0758_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 14352 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0759_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 16652 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _0760_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 15180 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0761_
timestamp 1723858470
transform 1 0 16100 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0762_
timestamp 1723858470
transform 1 0 16560 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0763_
timestamp 1723858470
transform 1 0 17572 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0764_
timestamp 1723858470
transform -1 0 18584 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0765_
timestamp 1723858470
transform 1 0 18400 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0766_
timestamp 1723858470
transform -1 0 19320 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _0767_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 17572 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0768_
timestamp 1723858470
transform 1 0 17756 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0769_
timestamp 1723858470
transform -1 0 18308 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0770_
timestamp 1723858470
transform 1 0 18400 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0771_
timestamp 1723858470
transform 1 0 18676 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1723858470
transform -1 0 18584 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0773_
timestamp 1723858470
transform 1 0 18676 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0774_
timestamp 1723858470
transform -1 0 19504 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0775_
timestamp 1723858470
transform -1 0 18400 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0776_
timestamp 1723858470
transform 1 0 18676 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0777_
timestamp 1723858470
transform -1 0 18768 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0778_
timestamp 1723858470
transform 1 0 18676 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0779_
timestamp 1723858470
transform -1 0 18768 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0780_
timestamp 1723858470
transform 1 0 20976 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0781_
timestamp 1723858470
transform -1 0 21988 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0782_
timestamp 1723858470
transform 1 0 20516 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0783_
timestamp 1723858470
transform 1 0 22356 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0784_
timestamp 1723858470
transform -1 0 22172 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0785_
timestamp 1723858470
transform 1 0 21528 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0786_
timestamp 1723858470
transform 1 0 22080 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0787_
timestamp 1723858470
transform -1 0 19688 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _0788_
timestamp 1723858470
transform 1 0 20516 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0789_
timestamp 1723858470
transform -1 0 20792 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1723858470
transform -1 0 20516 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o311ai_2  _0791_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 17388 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0792_
timestamp 1723858470
transform 1 0 18676 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0793_
timestamp 1723858470
transform -1 0 19044 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0794_
timestamp 1723858470
transform -1 0 20240 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0795_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 20608 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0796_
timestamp 1723858470
transform -1 0 20792 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0797_
timestamp 1723858470
transform 1 0 19964 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0798_
timestamp 1723858470
transform -1 0 21620 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0799_
timestamp 1723858470
transform -1 0 21528 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0800_
timestamp 1723858470
transform 1 0 21252 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _0801_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 22356 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0802_
timestamp 1723858470
transform -1 0 22448 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0803_
timestamp 1723858470
transform -1 0 21068 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0804_
timestamp 1723858470
transform 1 0 21068 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0805_
timestamp 1723858470
transform 1 0 22632 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0806_
timestamp 1723858470
transform 1 0 21252 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0807_
timestamp 1723858470
transform 1 0 21252 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0808_
timestamp 1723858470
transform 1 0 21252 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0809_
timestamp 1723858470
transform -1 0 21160 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0810_
timestamp 1723858470
transform 1 0 21988 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0811_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 21344 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0812_
timestamp 1723858470
transform 1 0 21712 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0813_
timestamp 1723858470
transform 1 0 22356 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0814_
timestamp 1723858470
transform 1 0 21252 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0815_
timestamp 1723858470
transform 1 0 22264 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0816_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 21160 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0817_
timestamp 1723858470
transform 1 0 21252 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0818_
timestamp 1723858470
transform 1 0 21896 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0819_
timestamp 1723858470
transform -1 0 22540 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0820_
timestamp 1723858470
transform -1 0 21896 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0821_
timestamp 1723858470
transform 1 0 21252 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0822_
timestamp 1723858470
transform 1 0 20792 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0823_
timestamp 1723858470
transform 1 0 20056 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0824_
timestamp 1723858470
transform -1 0 20792 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0825_
timestamp 1723858470
transform -1 0 20148 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1723858470
transform -1 0 19964 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0827_
timestamp 1723858470
transform 1 0 19688 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0828_
timestamp 1723858470
transform -1 0 19044 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0829_
timestamp 1723858470
transform 1 0 18400 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0830_
timestamp 1723858470
transform -1 0 17940 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0831_
timestamp 1723858470
transform -1 0 19504 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0832_
timestamp 1723858470
transform 1 0 17388 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0833_
timestamp 1723858470
transform 1 0 18676 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0834_
timestamp 1723858470
transform 1 0 16652 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0835_
timestamp 1723858470
transform 1 0 17572 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0836_
timestamp 1723858470
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1723858470
transform 1 0 17756 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0838_
timestamp 1723858470
transform 1 0 16284 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0839_
timestamp 1723858470
transform 1 0 16836 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0840_
timestamp 1723858470
transform 1 0 14996 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0841_
timestamp 1723858470
transform 1 0 16376 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0842_
timestamp 1723858470
transform -1 0 16008 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0843_
timestamp 1723858470
transform 1 0 14444 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0844_
timestamp 1723858470
transform 1 0 14996 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0845_
timestamp 1723858470
transform 1 0 14536 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0846_
timestamp 1723858470
transform 1 0 15088 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0847_
timestamp 1723858470
transform 1 0 14352 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0848_
timestamp 1723858470
transform 1 0 12236 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0849_
timestamp 1723858470
transform 1 0 13524 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0850_
timestamp 1723858470
transform 1 0 13616 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0851_
timestamp 1723858470
transform 1 0 11592 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0852_
timestamp 1723858470
transform 1 0 11868 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0853_
timestamp 1723858470
transform -1 0 12512 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0854_
timestamp 1723858470
transform -1 0 11592 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0855_
timestamp 1723858470
transform 1 0 11500 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0856_
timestamp 1723858470
transform 1 0 9752 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0857_
timestamp 1723858470
transform 1 0 10764 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0858_
timestamp 1723858470
transform 1 0 8464 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0859_
timestamp 1723858470
transform 1 0 9292 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0860_
timestamp 1723858470
transform 1 0 10396 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0861_
timestamp 1723858470
transform 1 0 8372 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0862_
timestamp 1723858470
transform 1 0 8556 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0863_
timestamp 1723858470
transform 1 0 7084 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0864_
timestamp 1723858470
transform -1 0 8648 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0865_
timestamp 1723858470
transform -1 0 7728 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0866_
timestamp 1723858470
transform 1 0 5336 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0867_
timestamp 1723858470
transform 1 0 6440 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0868_
timestamp 1723858470
transform 1 0 6900 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0869_
timestamp 1723858470
transform -1 0 6440 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0870_
timestamp 1723858470
transform 1 0 5796 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0871_
timestamp 1723858470
transform 1 0 7268 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0872_
timestamp 1723858470
transform -1 0 4600 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0873_
timestamp 1723858470
transform -1 0 7360 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1723858470
transform -1 0 5244 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 1723858470
transform -1 0 7360 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0876_
timestamp 1723858470
transform 1 0 5244 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0877_
timestamp 1723858470
transform 1 0 6348 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0878_
timestamp 1723858470
transform 1 0 7728 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0879_
timestamp 1723858470
transform 1 0 9384 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0880_
timestamp 1723858470
transform 1 0 12144 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0881_
timestamp 1723858470
transform 1 0 14996 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0882_
timestamp 1723858470
transform 1 0 17020 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0883_
timestamp 1723858470
transform 1 0 18768 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0884_
timestamp 1723858470
transform 1 0 20516 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0885_
timestamp 1723858470
transform -1 0 22448 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0886_
timestamp 1723858470
transform -1 0 22816 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0887_
timestamp 1723858470
transform 1 0 21528 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0888_
timestamp 1723858470
transform 1 0 22172 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0889_
timestamp 1723858470
transform -1 0 5704 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0890_
timestamp 1723858470
transform 1 0 5704 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0891_
timestamp 1723858470
transform -1 0 7820 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1723858470
transform 1 0 6440 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0893_
timestamp 1723858470
transform 1 0 4692 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0894_
timestamp 1723858470
transform 1 0 5796 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0895_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4600 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0896_
timestamp 1723858470
transform -1 0 4876 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0897_
timestamp 1723858470
transform -1 0 5704 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0898_
timestamp 1723858470
transform 1 0 4416 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0899_
timestamp 1723858470
transform 1 0 3956 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0900_
timestamp 1723858470
transform 1 0 5796 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0901_
timestamp 1723858470
transform 1 0 4416 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0902_
timestamp 1723858470
transform 1 0 5060 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0903_
timestamp 1723858470
transform 1 0 6348 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0904_
timestamp 1723858470
transform 1 0 6348 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0905_
timestamp 1723858470
transform 1 0 7544 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0906_
timestamp 1723858470
transform -1 0 8004 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0907_
timestamp 1723858470
transform 1 0 6900 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0908_
timestamp 1723858470
transform 1 0 7820 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 1723858470
transform -1 0 10028 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0910_
timestamp 1723858470
transform 1 0 8372 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0911_
timestamp 1723858470
transform 1 0 8832 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1723858470
transform 1 0 9016 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0913_
timestamp 1723858470
transform -1 0 9936 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0914_
timestamp 1723858470
transform 1 0 10120 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1723858470
transform -1 0 10856 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0916_
timestamp 1723858470
transform -1 0 10856 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0917_
timestamp 1723858470
transform -1 0 11408 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0918_
timestamp 1723858470
transform 1 0 10304 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0919_
timestamp 1723858470
transform -1 0 10764 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0920_
timestamp 1723858470
transform 1 0 11408 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0921_
timestamp 1723858470
transform 1 0 12052 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0922_
timestamp 1723858470
transform 1 0 10764 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1723858470
transform 1 0 13524 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0924_
timestamp 1723858470
transform -1 0 13892 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0925_
timestamp 1723858470
transform 1 0 12972 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0926_
timestamp 1723858470
transform 1 0 14168 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0927_
timestamp 1723858470
transform 1 0 14076 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0928_
timestamp 1723858470
transform -1 0 14536 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0929_
timestamp 1723858470
transform 1 0 14536 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0930_
timestamp 1723858470
transform 1 0 15180 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0931_
timestamp 1723858470
transform 1 0 14904 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0932_
timestamp 1723858470
transform 1 0 16652 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0933_
timestamp 1723858470
transform 1 0 16744 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0934_
timestamp 1723858470
transform 1 0 17204 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0935_
timestamp 1723858470
transform -1 0 18032 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0936_
timestamp 1723858470
transform -1 0 16836 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0937_
timestamp 1723858470
transform 1 0 16928 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0938_
timestamp 1723858470
transform 1 0 17480 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0939_
timestamp 1723858470
transform 1 0 16652 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0940_
timestamp 1723858470
transform -1 0 18768 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0941_
timestamp 1723858470
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0942_
timestamp 1723858470
transform -1 0 17664 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0943_
timestamp 1723858470
transform 1 0 17848 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1723858470
transform 1 0 18308 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0945_
timestamp 1723858470
transform 1 0 18676 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0946_
timestamp 1723858470
transform -1 0 18584 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0947_
timestamp 1723858470
transform -1 0 21068 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1723858470
transform -1 0 20332 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0949_
timestamp 1723858470
transform -1 0 20332 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0950_
timestamp 1723858470
transform -1 0 20792 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0951_
timestamp 1723858470
transform -1 0 20516 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0952_
timestamp 1723858470
transform 1 0 19228 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0953_
timestamp 1723858470
transform 1 0 21252 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0954_
timestamp 1723858470
transform -1 0 20976 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0955_
timestamp 1723858470
transform -1 0 21712 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0956_
timestamp 1723858470
transform 1 0 21160 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0957_
timestamp 1723858470
transform 1 0 22356 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0958_
timestamp 1723858470
transform -1 0 22356 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0959_
timestamp 1723858470
transform 1 0 21712 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0960_
timestamp 1723858470
transform -1 0 22632 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0961_
timestamp 1723858470
transform -1 0 22172 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0962_
timestamp 1723858470
transform -1 0 22356 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0963_
timestamp 1723858470
transform 1 0 22540 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0964_
timestamp 1723858470
transform -1 0 22540 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0965_
timestamp 1723858470
transform -1 0 21252 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0966_
timestamp 1723858470
transform -1 0 22724 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0967_
timestamp 1723858470
transform -1 0 21896 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0968_
timestamp 1723858470
transform -1 0 21344 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0969_
timestamp 1723858470
transform -1 0 21712 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0970_
timestamp 1723858470
transform 1 0 20424 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0971_
timestamp 1723858470
transform -1 0 21068 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0972_
timestamp 1723858470
transform -1 0 20792 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1723858470
transform -1 0 20148 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0974_
timestamp 1723858470
transform -1 0 19964 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0975_
timestamp 1723858470
transform -1 0 19688 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0976_
timestamp 1723858470
transform -1 0 19688 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0977_
timestamp 1723858470
transform -1 0 19044 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1723858470
transform 1 0 18216 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0979_
timestamp 1723858470
transform -1 0 21988 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0980_
timestamp 1723858470
transform -1 0 21620 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0981_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6348 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1723858470
transform 1 0 5796 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1723858470
transform -1 0 5704 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1723858470
transform -1 0 7176 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1723858470
transform 1 0 6992 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1723858470
transform 1 0 8556 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1723858470
transform 1 0 8832 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1723858470
transform 1 0 10948 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1723858470
transform 1 0 11316 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1723858470
transform -1 0 13432 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1723858470
transform 1 0 13892 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1723858470
transform 1 0 14076 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1723858470
transform 1 0 14628 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1723858470
transform 1 0 15456 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1723858470
transform 1 0 16100 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1723858470
transform 1 0 16468 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1723858470
transform 1 0 18676 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1723858470
transform 1 0 18768 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1723858470
transform 1 0 19504 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1723858470
transform 1 0 20792 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1723858470
transform -1 0 22816 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1723858470
transform 1 0 21252 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1723858470
transform -1 0 5704 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1723858470
transform -1 0 6900 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1723858470
transform 1 0 5796 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1723858470
transform 1 0 5244 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1723858470
transform 1 0 4876 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1723858470
transform 1 0 4876 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1723858470
transform -1 0 7268 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1723858470
transform 1 0 7360 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1723858470
transform -1 0 9292 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1723858470
transform 1 0 8556 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1723858470
transform 1 0 10212 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1723858470
transform 1 0 10948 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1723858470
transform 1 0 11408 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1723858470
transform 1 0 13340 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1723858470
transform 1 0 13800 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1723858470
transform -1 0 16744 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1723858470
transform -1 0 17940 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1723858470
transform -1 0 18308 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1723858470
transform -1 0 18584 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1723858470
transform 1 0 19136 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1723858470
transform 1 0 17664 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1723858470
transform 1 0 19596 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1723858470
transform 1 0 19688 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1723858470
transform 1 0 20332 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1723858470
transform 1 0 21620 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1723858470
transform 1 0 21620 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1723858470
transform 1 0 21528 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1723858470
transform 1 0 21344 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1723858470
transform 1 0 21252 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1723858470
transform 1 0 19780 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1723858470
transform 1 0 18860 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1723858470
transform 1 0 18676 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1723858470
transform 1 0 21620 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  fanout11 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 10304 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout12
timestamp 1723858470
transform -1 0 19596 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout13
timestamp 1723858470
transform 1 0 21252 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout14
timestamp 1723858470
transform -1 0 23000 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout15 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 20700 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout16 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21620 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout17 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 17572 0 1 22304
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp 1723858470
transform -1 0 6256 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 1723858470
transform -1 0 5520 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1723858470
transform 1 0 6256 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1723858470
transform 1 0 22172 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1723858470
transform -1 0 22816 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout23
timestamp 1723858470
transform -1 0 9016 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout24
timestamp 1723858470
transform 1 0 12972 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1723858470
transform -1 0 13432 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1723858470
transform -1 0 16468 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1723858470
transform 1 0 20792 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1723858470
transform 1 0 20424 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp 1723858470
transform -1 0 23092 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1723858470
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1723858470
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1723858470
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1723858470
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1723858470
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1723858470
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1723858470
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1723858470
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1723858470
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1723858470
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1723858470
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1723858470
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1723858470
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1723858470
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1723858470
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1723858470
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1723858470
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1723858470
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1723858470
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1723858470
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1723858470
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1723858470
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_237 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 22356 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1723858470
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1723858470
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1723858470
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1723858470
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1723858470
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1723858470
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1723858470
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1723858470
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1723858470
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1723858470
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1723858470
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1723858470
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1723858470
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1723858470
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1723858470
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1723858470
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1723858470
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1723858470
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1723858470
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1723858470
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1723858470
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1723858470
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1723858470
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_237
timestamp 1723858470
transform 1 0 22356 0 -1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1723858470
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1723858470
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1723858470
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1723858470
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1723858470
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1723858470
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1723858470
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1723858470
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1723858470
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1723858470
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1723858470
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1723858470
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1723858470
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1723858470
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1723858470
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1723858470
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1723858470
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1723858470
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1723858470
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1723858470
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1723858470
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1723858470
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1723858470
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1723858470
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1723858470
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1723858470
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1723858470
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1723858470
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1723858470
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1723858470
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1723858470
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1723858470
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1723858470
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1723858470
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1723858470
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1723858470
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1723858470
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1723858470
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1723858470
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1723858470
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1723858470
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1723858470
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1723858470
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1723858470
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1723858470
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1723858470
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1723858470
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1723858470
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1723858470
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1723858470
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_237
timestamp 1723858470
transform 1 0 22356 0 -1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1723858470
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1723858470
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1723858470
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1723858470
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1723858470
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1723858470
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1723858470
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1723858470
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1723858470
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1723858470
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1723858470
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1723858470
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1723858470
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1723858470
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1723858470
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1723858470
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1723858470
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1723858470
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1723858470
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1723858470
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1723858470
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1723858470
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1723858470
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1723858470
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1723858470
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1723858470
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1723858470
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1723858470
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1723858470
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1723858470
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1723858470
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1723858470
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1723858470
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1723858470
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1723858470
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1723858470
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1723858470
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1723858470
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1723858470
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1723858470
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1723858470
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1723858470
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1723858470
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1723858470
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1723858470
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1723858470
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1723858470
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1723858470
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1723858470
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1723858470
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_237
timestamp 1723858470
transform 1 0 22356 0 -1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1723858470
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1723858470
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1723858470
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1723858470
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1723858470
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1723858470
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1723858470
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1723858470
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1723858470
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1723858470
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1723858470
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1723858470
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1723858470
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1723858470
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1723858470
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1723858470
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1723858470
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1723858470
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1723858470
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1723858470
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1723858470
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1723858470
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1723858470
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1723858470
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_233
timestamp 1723858470
transform 1 0 21988 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_241
timestamp 1723858470
transform 1 0 22724 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1723858470
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1723858470
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1723858470
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1723858470
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1723858470
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1723858470
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1723858470
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1723858470
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1723858470
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1723858470
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1723858470
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1723858470
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1723858470
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1723858470
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1723858470
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1723858470
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1723858470
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1723858470
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1723858470
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1723858470
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1723858470
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1723858470
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1723858470
transform 1 0 20516 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1723858470
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1723858470
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_237
timestamp 1723858470
transform 1 0 22356 0 -1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1723858470
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1723858470
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1723858470
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1723858470
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1723858470
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1723858470
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1723858470
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1723858470
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1723858470
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1723858470
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1723858470
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1723858470
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1723858470
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1723858470
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1723858470
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1723858470
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1723858470
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1723858470
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1723858470
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1723858470
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1723858470
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1723858470
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1723858470
transform 1 0 19780 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1723858470
transform 1 0 20884 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1723858470
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1723858470
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1723858470
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1723858470
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1723858470
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1723858470
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1723858470
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1723858470
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1723858470
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1723858470
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1723858470
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1723858470
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1723858470
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1723858470
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1723858470
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1723858470
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1723858470
transform 1 0 14260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1723858470
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1723858470
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1723858470
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1723858470
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1723858470
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1723858470
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1723858470
transform 1 0 20516 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1723858470
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1723858470
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_237
timestamp 1723858470
transform 1 0 22356 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1723858470
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1723858470
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1723858470
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1723858470
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1723858470
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_69
timestamp 1723858470
transform 1 0 6900 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1723858470
transform 1 0 8004 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1723858470
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1723858470
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1723858470
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1723858470
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1723858470
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1723858470
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1723858470
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1723858470
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1723858470
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1723858470
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1723858470
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1723858470
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1723858470
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1723858470
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1723858470
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1723858470
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1723858470
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1723858470
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1723858470
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_39
timestamp 1723858470
transform 1 0 4140 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_76
timestamp 1723858470
transform 1 0 7544 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_88
timestamp 1723858470
transform 1 0 8648 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_100
timestamp 1723858470
transform 1 0 9752 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_106
timestamp 1723858470
transform 1 0 10304 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1723858470
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1723858470
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1723858470
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1723858470
transform 1 0 14260 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1723858470
transform 1 0 15364 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1723858470
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1723858470
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1723858470
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1723858470
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1723858470
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1723858470
transform 1 0 20516 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1723858470
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1723858470
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_237
timestamp 1723858470
transform 1 0 22356 0 -1 7072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1723858470
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1723858470
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1723858470
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1723858470
transform 1 0 3220 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_37
timestamp 1723858470
transform 1 0 3956 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_79
timestamp 1723858470
transform 1 0 7820 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1723858470
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_85
timestamp 1723858470
transform 1 0 8372 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_92
timestamp 1723858470
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_104
timestamp 1723858470
transform 1 0 10120 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1723858470
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1723858470
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1723858470
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_141
timestamp 1723858470
transform 1 0 13524 0 1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1723858470
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1723858470
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1723858470
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1723858470
transform 1 0 17940 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1723858470
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1723858470
transform 1 0 18676 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1723858470
transform 1 0 19780 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_221 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_226
timestamp 1723858470
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_238
timestamp 1723858470
transform 1 0 22448 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_244
timestamp 1723858470
transform 1 0 23000 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1723858470
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1723858470
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1723858470
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_39
timestamp 1723858470
transform 1 0 4140 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_70
timestamp 1723858470
transform 1 0 6992 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_78
timestamp 1723858470
transform 1 0 7728 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_129
timestamp 1723858470
transform 1 0 12420 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_155
timestamp 1723858470
transform 1 0 14812 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_163
timestamp 1723858470
transform 1 0 15548 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1723858470
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1723858470
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1723858470
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_193
timestamp 1723858470
transform 1 0 18308 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_201
timestamp 1723858470
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_213
timestamp 1723858470
transform 1 0 20148 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_217
timestamp 1723858470
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1723858470
transform 1 0 21068 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_241
timestamp 1723858470
transform 1 0 22724 0 -1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1723858470
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1723858470
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1723858470
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1723858470
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1723858470
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_53
timestamp 1723858470
transform 1 0 5428 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_61
timestamp 1723858470
transform 1 0 6164 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_73
timestamp 1723858470
transform 1 0 7268 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1723858470
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_103
timestamp 1723858470
transform 1 0 10028 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_134
timestamp 1723858470
transform 1 0 12880 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_186
timestamp 1723858470
transform 1 0 17664 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1723858470
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_197
timestamp 1723858470
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_215
timestamp 1723858470
transform 1 0 20332 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1723858470
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1723858470
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1723858470
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1723858470
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1723858470
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_103
timestamp 1723858470
transform 1 0 10028 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_130
timestamp 1723858470
transform 1 0 12512 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_164
timestamp 1723858470
transform 1 0 15640 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_189
timestamp 1723858470
transform 1 0 17940 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_225
timestamp 1723858470
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_242
timestamp 1723858470
transform 1 0 22816 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1723858470
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1723858470
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1723858470
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1723858470
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_41
timestamp 1723858470
transform 1 0 4324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_70
timestamp 1723858470
transform 1 0 6992 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1723858470
transform 1 0 8004 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1723858470
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_109
timestamp 1723858470
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_118
timestamp 1723858470
transform 1 0 11408 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_122
timestamp 1723858470
transform 1 0 11776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_130
timestamp 1723858470
transform 1 0 12512 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1723858470
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_141
timestamp 1723858470
transform 1 0 13524 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_147
timestamp 1723858470
transform 1 0 14076 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_153
timestamp 1723858470
transform 1 0 14628 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_163
timestamp 1723858470
transform 1 0 15548 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_190
timestamp 1723858470
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_197
timestamp 1723858470
transform 1 0 18676 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_208
timestamp 1723858470
transform 1 0 19688 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_225
timestamp 1723858470
transform 1 0 21252 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_244
timestamp 1723858470
transform 1 0 23000 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1723858470
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1723858470
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_27
timestamp 1723858470
transform 1 0 3036 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_35
timestamp 1723858470
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_73
timestamp 1723858470
transform 1 0 7268 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_85
timestamp 1723858470
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_94
timestamp 1723858470
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_102
timestamp 1723858470
transform 1 0 9936 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_110
timestamp 1723858470
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_113
timestamp 1723858470
transform 1 0 10948 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_132
timestamp 1723858470
transform 1 0 12696 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_140
timestamp 1723858470
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_149
timestamp 1723858470
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_164
timestamp 1723858470
transform 1 0 15640 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_169
timestamp 1723858470
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1723858470
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_205
timestamp 1723858470
transform 1 0 19412 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_211
timestamp 1723858470
transform 1 0 19964 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_244
timestamp 1723858470
transform 1 0 23000 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1723858470
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1723858470
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1723858470
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1723858470
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_41
timestamp 1723858470
transform 1 0 4324 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_68
timestamp 1723858470
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_80
timestamp 1723858470
transform 1 0 7912 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_92
timestamp 1723858470
transform 1 0 9016 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_111
timestamp 1723858470
transform 1 0 10764 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1723858470
transform 1 0 12788 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1723858470
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_144
timestamp 1723858470
transform 1 0 13800 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_150
timestamp 1723858470
transform 1 0 14352 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_161
timestamp 1723858470
transform 1 0 15364 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_173
timestamp 1723858470
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1723858470
transform 1 0 18676 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_209
timestamp 1723858470
transform 1 0 19780 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_217
timestamp 1723858470
transform 1 0 20516 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_242
timestamp 1723858470
transform 1 0 22816 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1723858470
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1723858470
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1723858470
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_39
timestamp 1723858470
transform 1 0 4140 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_45
timestamp 1723858470
transform 1 0 4692 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_88
timestamp 1723858470
transform 1 0 8648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1723858470
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1723858470
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_163
timestamp 1723858470
transform 1 0 15548 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1723858470
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_198
timestamp 1723858470
transform 1 0 18768 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_210
timestamp 1723858470
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_220
timestamp 1723858470
transform 1 0 20792 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_225
timestamp 1723858470
transform 1 0 21252 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_240
timestamp 1723858470
transform 1 0 22632 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_244
timestamp 1723858470
transform 1 0 23000 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1723858470
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1723858470
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1723858470
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1723858470
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1723858470
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_53
timestamp 1723858470
transform 1 0 5428 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_73
timestamp 1723858470
transform 1 0 7268 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 1723858470
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1723858470
transform 1 0 8372 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_106
timestamp 1723858470
transform 1 0 10304 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_112
timestamp 1723858470
transform 1 0 10856 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_129
timestamp 1723858470
transform 1 0 12420 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1723858470
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1723858470
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_176
timestamp 1723858470
transform 1 0 16744 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_185
timestamp 1723858470
transform 1 0 17572 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_193
timestamp 1723858470
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_197
timestamp 1723858470
transform 1 0 18676 0 1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1723858470
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1723858470
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1723858470
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1723858470
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_51
timestamp 1723858470
transform 1 0 5244 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_74
timestamp 1723858470
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_86
timestamp 1723858470
transform 1 0 8464 0 -1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_99
timestamp 1723858470
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1723858470
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 1723858470
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_133
timestamp 1723858470
transform 1 0 12788 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_163
timestamp 1723858470
transform 1 0 15548 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1723858470
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_169
timestamp 1723858470
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_178
timestamp 1723858470
transform 1 0 16928 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1723858470
transform 1 0 21068 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1723858470
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1723858470
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1723858470
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1723858470
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_41
timestamp 1723858470
transform 1 0 4324 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_68
timestamp 1723858470
transform 1 0 6808 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_74
timestamp 1723858470
transform 1 0 7360 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1723858470
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_103
timestamp 1723858470
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_112
timestamp 1723858470
transform 1 0 10856 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_118
timestamp 1723858470
transform 1 0 11408 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_141
timestamp 1723858470
transform 1 0 13524 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_170
timestamp 1723858470
transform 1 0 16192 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_182
timestamp 1723858470
transform 1 0 17296 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1723858470
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1723858470
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1723858470
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1723858470
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1723858470
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1723858470
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_66
timestamp 1723858470
transform 1 0 6624 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_86
timestamp 1723858470
transform 1 0 8464 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_108
timestamp 1723858470
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_113
timestamp 1723858470
transform 1 0 10948 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_119
timestamp 1723858470
transform 1 0 11500 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_127
timestamp 1723858470
transform 1 0 12236 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_135
timestamp 1723858470
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_159
timestamp 1723858470
transform 1 0 15180 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1723858470
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_178
timestamp 1723858470
transform 1 0 16928 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_190
timestamp 1723858470
transform 1 0 18032 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_198
timestamp 1723858470
transform 1 0 18768 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_206
timestamp 1723858470
transform 1 0 19504 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1723858470
transform 1 0 20976 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_244
timestamp 1723858470
transform 1 0 23000 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1723858470
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1723858470
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1723858470
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1723858470
transform 1 0 3220 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_37
timestamp 1723858470
transform 1 0 3956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1723858470
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_85
timestamp 1723858470
transform 1 0 8372 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_95
timestamp 1723858470
transform 1 0 9292 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_106
timestamp 1723858470
transform 1 0 10304 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_115
timestamp 1723858470
transform 1 0 11132 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_127
timestamp 1723858470
transform 1 0 12236 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_141
timestamp 1723858470
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_148
timestamp 1723858470
transform 1 0 14168 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_156
timestamp 1723858470
transform 1 0 14904 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_183
timestamp 1723858470
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1723858470
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_197
timestamp 1723858470
transform 1 0 18676 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_204
timestamp 1723858470
transform 1 0 19320 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_231
timestamp 1723858470
transform 1 0 21804 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_236
timestamp 1723858470
transform 1 0 22264 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_244
timestamp 1723858470
transform 1 0 23000 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1723858470
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1723858470
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1723858470
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1723858470
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1723858470
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1723858470
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_66
timestamp 1723858470
transform 1 0 6624 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_78
timestamp 1723858470
transform 1 0 7728 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_90
timestamp 1723858470
transform 1 0 8832 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1723858470
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_125
timestamp 1723858470
transform 1 0 12052 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_142
timestamp 1723858470
transform 1 0 13616 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_159
timestamp 1723858470
transform 1 0 15180 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1723858470
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_169
timestamp 1723858470
transform 1 0 16100 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_179
timestamp 1723858470
transform 1 0 17020 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_192
timestamp 1723858470
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_206
timestamp 1723858470
transform 1 0 19504 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_218
timestamp 1723858470
transform 1 0 20608 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_225
timestamp 1723858470
transform 1 0 21252 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_244
timestamp 1723858470
transform 1 0 23000 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1723858470
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1723858470
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1723858470
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1723858470
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1723858470
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1723858470
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1723858470
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1723858470
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1723858470
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_85
timestamp 1723858470
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_100
timestamp 1723858470
transform 1 0 9752 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_104
timestamp 1723858470
transform 1 0 10120 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_110
timestamp 1723858470
transform 1 0 10672 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_116
timestamp 1723858470
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_129
timestamp 1723858470
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 1723858470
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_157
timestamp 1723858470
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_169
timestamp 1723858470
transform 1 0 16100 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_194
timestamp 1723858470
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_202
timestamp 1723858470
transform 1 0 19136 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_215
timestamp 1723858470
transform 1 0 20332 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_220
timestamp 1723858470
transform 1 0 20792 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_224
timestamp 1723858470
transform 1 0 21160 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_242
timestamp 1723858470
transform 1 0 22816 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1723858470
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1723858470
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1723858470
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_39
timestamp 1723858470
transform 1 0 4140 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_47
timestamp 1723858470
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_73
timestamp 1723858470
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_79
timestamp 1723858470
transform 1 0 7820 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_92
timestamp 1723858470
transform 1 0 9016 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_103
timestamp 1723858470
transform 1 0 10028 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1723858470
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_113
timestamp 1723858470
transform 1 0 10948 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_128
timestamp 1723858470
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_136
timestamp 1723858470
transform 1 0 13064 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_142
timestamp 1723858470
transform 1 0 13616 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_156
timestamp 1723858470
transform 1 0 14904 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_185
timestamp 1723858470
transform 1 0 17572 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_189
timestamp 1723858470
transform 1 0 17940 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_193
timestamp 1723858470
transform 1 0 18308 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_201
timestamp 1723858470
transform 1 0 19044 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_207
timestamp 1723858470
transform 1 0 19596 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_211
timestamp 1723858470
transform 1 0 19964 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1723858470
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_239
timestamp 1723858470
transform 1 0 22540 0 -1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1723858470
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1723858470
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1723858470
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1723858470
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_41
timestamp 1723858470
transform 1 0 4324 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_51
timestamp 1723858470
transform 1 0 5244 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_59
timestamp 1723858470
transform 1 0 5980 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_92
timestamp 1723858470
transform 1 0 9016 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_102
timestamp 1723858470
transform 1 0 9936 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_110
timestamp 1723858470
transform 1 0 10672 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_116
timestamp 1723858470
transform 1 0 11224 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_120
timestamp 1723858470
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_145
timestamp 1723858470
transform 1 0 13892 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_164
timestamp 1723858470
transform 1 0 15640 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_168
timestamp 1723858470
transform 1 0 16008 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_183
timestamp 1723858470
transform 1 0 17388 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1723858470
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_197
timestamp 1723858470
transform 1 0 18676 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_203
timestamp 1723858470
transform 1 0 19228 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_213
timestamp 1723858470
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_223
timestamp 1723858470
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_240
timestamp 1723858470
transform 1 0 22632 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_244
timestamp 1723858470
transform 1 0 23000 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1723858470
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1723858470
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1723858470
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_39
timestamp 1723858470
transform 1 0 4140 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_50
timestamp 1723858470
transform 1 0 5152 0 -1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_77
timestamp 1723858470
transform 1 0 7636 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_89
timestamp 1723858470
transform 1 0 8740 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_106
timestamp 1723858470
transform 1 0 10304 0 -1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1723858470
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1723858470
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1723858470
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_149
timestamp 1723858470
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_160
timestamp 1723858470
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_183
timestamp 1723858470
transform 1 0 17388 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_191
timestamp 1723858470
transform 1 0 18124 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_197
timestamp 1723858470
transform 1 0 18676 0 -1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_204
timestamp 1723858470
transform 1 0 19320 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_216
timestamp 1723858470
transform 1 0 20424 0 -1 16864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_231
timestamp 1723858470
transform 1 0 21804 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_243
timestamp 1723858470
transform 1 0 22908 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1723858470
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1723858470
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1723858470
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1723858470
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_41
timestamp 1723858470
transform 1 0 4324 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_67
timestamp 1723858470
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_71
timestamp 1723858470
transform 1 0 7084 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1723858470
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_85
timestamp 1723858470
transform 1 0 8372 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_89
timestamp 1723858470
transform 1 0 8740 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_116
timestamp 1723858470
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_128
timestamp 1723858470
transform 1 0 12328 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_141
timestamp 1723858470
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_158
timestamp 1723858470
transform 1 0 15088 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_165
timestamp 1723858470
transform 1 0 15732 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_190
timestamp 1723858470
transform 1 0 18032 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_213
timestamp 1723858470
transform 1 0 20148 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_242
timestamp 1723858470
transform 1 0 22816 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1723858470
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1723858470
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1723858470
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_39
timestamp 1723858470
transform 1 0 4140 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_43
timestamp 1723858470
transform 1 0 4508 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_64
timestamp 1723858470
transform 1 0 6440 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_78
timestamp 1723858470
transform 1 0 7728 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_89
timestamp 1723858470
transform 1 0 8740 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_97
timestamp 1723858470
transform 1 0 9476 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_107
timestamp 1723858470
transform 1 0 10396 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1723858470
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_116
timestamp 1723858470
transform 1 0 11224 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_120
timestamp 1723858470
transform 1 0 11592 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1723858470
transform 1 0 14260 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_161
timestamp 1723858470
transform 1 0 15364 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_182
timestamp 1723858470
transform 1 0 17296 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_214
timestamp 1723858470
transform 1 0 20240 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 1723858470
transform 1 0 20976 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_225
timestamp 1723858470
transform 1 0 21252 0 -1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1723858470
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1723858470
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1723858470
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1723858470
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1723858470
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_90
timestamp 1723858470
transform 1 0 8832 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_101
timestamp 1723858470
transform 1 0 9844 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_108
timestamp 1723858470
transform 1 0 10488 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_118
timestamp 1723858470
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_130
timestamp 1723858470
transform 1 0 12512 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1723858470
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_141
timestamp 1723858470
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_149
timestamp 1723858470
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_164
timestamp 1723858470
transform 1 0 15640 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_168
timestamp 1723858470
transform 1 0 16008 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_179
timestamp 1723858470
transform 1 0 17020 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_204
timestamp 1723858470
transform 1 0 19320 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_212
timestamp 1723858470
transform 1 0 20056 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_220
timestamp 1723858470
transform 1 0 20792 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1723858470
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1723858470
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1723858470
transform 1 0 3036 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_39
timestamp 1723858470
transform 1 0 4140 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_47
timestamp 1723858470
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_65
timestamp 1723858470
transform 1 0 6532 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_85
timestamp 1723858470
transform 1 0 8372 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_106
timestamp 1723858470
transform 1 0 10304 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_133
timestamp 1723858470
transform 1 0 12788 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_141
timestamp 1723858470
transform 1 0 13524 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_146
timestamp 1723858470
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1723858470
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_176
timestamp 1723858470
transform 1 0 16744 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_188
timestamp 1723858470
transform 1 0 17848 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_201
timestamp 1723858470
transform 1 0 19044 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_205
timestamp 1723858470
transform 1 0 19412 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1723858470
transform 1 0 20976 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_244
timestamp 1723858470
transform 1 0 23000 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1723858470
transform 1 0 828 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1723858470
transform 1 0 1932 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1723858470
transform 1 0 3036 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1723858470
transform 1 0 3220 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1723858470
transform 1 0 4324 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_58
timestamp 1723858470
transform 1 0 5888 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_66
timestamp 1723858470
transform 1 0 6624 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_73
timestamp 1723858470
transform 1 0 7268 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_85
timestamp 1723858470
transform 1 0 8372 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_135
timestamp 1723858470
transform 1 0 12972 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1723858470
transform 1 0 13340 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_155
timestamp 1723858470
transform 1 0 14812 0 1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_175
timestamp 1723858470
transform 1 0 16652 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_187
timestamp 1723858470
transform 1 0 17756 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_200
timestamp 1723858470
transform 1 0 18952 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_208
timestamp 1723858470
transform 1 0 19688 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_242
timestamp 1723858470
transform 1 0 22816 0 1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1723858470
transform 1 0 828 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1723858470
transform 1 0 1932 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1723858470
transform 1 0 3036 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1723858470
transform 1 0 4140 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1723858470
transform 1 0 5244 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1723858470
transform 1 0 5612 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1723858470
transform 1 0 5796 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_62
timestamp 1723858470
transform 1 0 6256 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_71
timestamp 1723858470
transform 1 0 7084 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_80
timestamp 1723858470
transform 1 0 7912 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_113
timestamp 1723858470
transform 1 0 10948 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_122
timestamp 1723858470
transform 1 0 11776 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_126
timestamp 1723858470
transform 1 0 12144 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_134
timestamp 1723858470
transform 1 0 12880 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_153
timestamp 1723858470
transform 1 0 14628 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_165
timestamp 1723858470
transform 1 0 15732 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_169
timestamp 1723858470
transform 1 0 16100 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_177
timestamp 1723858470
transform 1 0 16836 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_188
timestamp 1723858470
transform 1 0 17848 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_206
timestamp 1723858470
transform 1 0 19504 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1723858470
transform 1 0 828 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1723858470
transform 1 0 1932 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1723858470
transform 1 0 3036 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1723858470
transform 1 0 3220 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_41
timestamp 1723858470
transform 1 0 4324 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_65
timestamp 1723858470
transform 1 0 6532 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_72
timestamp 1723858470
transform 1 0 7176 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_91
timestamp 1723858470
transform 1 0 8924 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_103
timestamp 1723858470
transform 1 0 10028 0 1 20128
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1723858470
transform 1 0 10580 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_121
timestamp 1723858470
transform 1 0 11684 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_129
timestamp 1723858470
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_136
timestamp 1723858470
transform 1 0 13064 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_146
timestamp 1723858470
transform 1 0 13984 0 1 20128
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_154
timestamp 1723858470
transform 1 0 14720 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_166
timestamp 1723858470
transform 1 0 15824 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_190
timestamp 1723858470
transform 1 0 18032 0 1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_200
timestamp 1723858470
transform 1 0 18952 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_212
timestamp 1723858470
transform 1 0 20056 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_228
timestamp 1723858470
transform 1 0 21528 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_239
timestamp 1723858470
transform 1 0 22540 0 1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1723858470
transform 1 0 828 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1723858470
transform 1 0 1932 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1723858470
transform 1 0 3036 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_39
timestamp 1723858470
transform 1 0 4140 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1723858470
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_69
timestamp 1723858470
transform 1 0 6900 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_92
timestamp 1723858470
transform 1 0 9016 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_101
timestamp 1723858470
transform 1 0 9844 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_107
timestamp 1723858470
transform 1 0 10396 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_113
timestamp 1723858470
transform 1 0 10948 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_121
timestamp 1723858470
transform 1 0 11684 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_133
timestamp 1723858470
transform 1 0 12788 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_141
timestamp 1723858470
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_148
timestamp 1723858470
transform 1 0 14168 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_164
timestamp 1723858470
transform 1 0 15640 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_169
timestamp 1723858470
transform 1 0 16100 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_174
timestamp 1723858470
transform 1 0 16560 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_180
timestamp 1723858470
transform 1 0 17112 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_184
timestamp 1723858470
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_196
timestamp 1723858470
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_208
timestamp 1723858470
transform 1 0 19688 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1723858470
transform 1 0 20976 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_238
timestamp 1723858470
transform 1 0 22448 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_244
timestamp 1723858470
transform 1 0 23000 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1723858470
transform 1 0 828 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1723858470
transform 1 0 1932 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1723858470
transform 1 0 3036 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1723858470
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_41
timestamp 1723858470
transform 1 0 4324 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_47
timestamp 1723858470
transform 1 0 4876 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_54
timestamp 1723858470
transform 1 0 5520 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1723858470
transform 1 0 8188 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_131
timestamp 1723858470
transform 1 0 12604 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_135
timestamp 1723858470
transform 1 0 12972 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_162
timestamp 1723858470
transform 1 0 15456 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_170
timestamp 1723858470
transform 1 0 16192 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_183
timestamp 1723858470
transform 1 0 17388 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_208
timestamp 1723858470
transform 1 0 19688 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_214
timestamp 1723858470
transform 1 0 20240 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_220
timestamp 1723858470
transform 1 0 20792 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_237
timestamp 1723858470
transform 1 0 22356 0 1 21216
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1723858470
transform 1 0 828 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1723858470
transform 1 0 1932 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1723858470
transform 1 0 3036 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_39
timestamp 1723858470
transform 1 0 4140 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_47
timestamp 1723858470
transform 1 0 4876 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_54
timestamp 1723858470
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_57
timestamp 1723858470
transform 1 0 5796 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_66
timestamp 1723858470
transform 1 0 6624 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1723858470
transform 1 0 10764 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_113
timestamp 1723858470
transform 1 0 10948 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_140
timestamp 1723858470
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_199
timestamp 1723858470
transform 1 0 18860 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1723858470
transform 1 0 21068 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_242
timestamp 1723858470
transform 1 0 22816 0 -1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1723858470
transform 1 0 828 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1723858470
transform 1 0 1932 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1723858470
transform 1 0 3036 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1723858470
transform 1 0 3220 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_41
timestamp 1723858470
transform 1 0 4324 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_88
timestamp 1723858470
transform 1 0 8648 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_97
timestamp 1723858470
transform 1 0 9476 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_108
timestamp 1723858470
transform 1 0 10488 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_127
timestamp 1723858470
transform 1 0 12236 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_134
timestamp 1723858470
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_157
timestamp 1723858470
transform 1 0 14996 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_190
timestamp 1723858470
transform 1 0 18032 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_215
timestamp 1723858470
transform 1 0 20332 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_235
timestamp 1723858470
transform 1 0 22172 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_243
timestamp 1723858470
transform 1 0 22908 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_3
timestamp 1723858470
transform 1 0 828 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_11
timestamp 1723858470
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_16
timestamp 1723858470
transform 1 0 2024 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_29
timestamp 1723858470
transform 1 0 3220 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_41
timestamp 1723858470
transform 1 0 4324 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_48
timestamp 1723858470
transform 1 0 4968 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_57
timestamp 1723858470
transform 1 0 5796 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_66
timestamp 1723858470
transform 1 0 6624 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_74
timestamp 1723858470
transform 1 0 7360 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_82
timestamp 1723858470
transform 1 0 8096 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_85
timestamp 1723858470
transform 1 0 8372 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_97
timestamp 1723858470
transform 1 0 9476 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_105
timestamp 1723858470
transform 1 0 10212 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_113
timestamp 1723858470
transform 1 0 10948 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_121
timestamp 1723858470
transform 1 0 11684 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_133
timestamp 1723858470
transform 1 0 12788 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_139
timestamp 1723858470
transform 1 0 13340 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_147
timestamp 1723858470
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_159
timestamp 1723858470
transform 1 0 15180 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1723858470
transform 1 0 15916 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_169
timestamp 1723858470
transform 1 0 16100 0 -1 23392
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_176
timestamp 1723858470
transform 1 0 16744 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_188
timestamp 1723858470
transform 1 0 17848 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_197
timestamp 1723858470
transform 1 0 18676 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_214
timestamp 1723858470
transform 1 0 20240 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_222
timestamp 1723858470
transform 1 0 20976 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_233
timestamp 1723858470
transform 1 0 21988 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_243
timestamp 1723858470
transform 1 0 22908 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 23092 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 22816 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1723858470
transform 1 0 1748 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1723858470
transform 1 0 4692 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1723858470
transform -1 0 8096 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1723858470
transform 1 0 10304 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 13524 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1723858470
transform 1 0 16468 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1723858470
transform 1 0 19412 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1723858470
transform 1 0 22356 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_42
timestamp 1723858470
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1723858470
transform -1 0 23368 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_43
timestamp 1723858470
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1723858470
transform -1 0 23368 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_44
timestamp 1723858470
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1723858470
transform -1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_45
timestamp 1723858470
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1723858470
transform -1 0 23368 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_46
timestamp 1723858470
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1723858470
transform -1 0 23368 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_47
timestamp 1723858470
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1723858470
transform -1 0 23368 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_48
timestamp 1723858470
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1723858470
transform -1 0 23368 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_49
timestamp 1723858470
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1723858470
transform -1 0 23368 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_50
timestamp 1723858470
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1723858470
transform -1 0 23368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_51
timestamp 1723858470
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1723858470
transform -1 0 23368 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_52
timestamp 1723858470
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1723858470
transform -1 0 23368 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_53
timestamp 1723858470
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1723858470
transform -1 0 23368 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_54
timestamp 1723858470
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1723858470
transform -1 0 23368 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_55
timestamp 1723858470
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1723858470
transform -1 0 23368 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_56
timestamp 1723858470
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1723858470
transform -1 0 23368 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_57
timestamp 1723858470
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1723858470
transform -1 0 23368 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_58
timestamp 1723858470
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1723858470
transform -1 0 23368 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_59
timestamp 1723858470
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1723858470
transform -1 0 23368 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_60
timestamp 1723858470
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1723858470
transform -1 0 23368 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_61
timestamp 1723858470
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1723858470
transform -1 0 23368 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_62
timestamp 1723858470
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1723858470
transform -1 0 23368 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_63
timestamp 1723858470
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1723858470
transform -1 0 23368 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_64
timestamp 1723858470
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1723858470
transform -1 0 23368 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_65
timestamp 1723858470
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1723858470
transform -1 0 23368 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_66
timestamp 1723858470
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1723858470
transform -1 0 23368 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_67
timestamp 1723858470
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1723858470
transform -1 0 23368 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_68
timestamp 1723858470
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1723858470
transform -1 0 23368 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_69
timestamp 1723858470
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1723858470
transform -1 0 23368 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_70
timestamp 1723858470
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1723858470
transform -1 0 23368 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_71
timestamp 1723858470
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1723858470
transform -1 0 23368 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_72
timestamp 1723858470
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1723858470
transform -1 0 23368 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_73
timestamp 1723858470
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1723858470
transform -1 0 23368 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_74
timestamp 1723858470
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1723858470
transform -1 0 23368 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_75
timestamp 1723858470
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1723858470
transform -1 0 23368 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_76
timestamp 1723858470
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1723858470
transform -1 0 23368 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_77
timestamp 1723858470
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1723858470
transform -1 0 23368 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_78
timestamp 1723858470
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1723858470
transform -1 0 23368 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_79
timestamp 1723858470
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1723858470
transform -1 0 23368 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_80
timestamp 1723858470
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1723858470
transform -1 0 23368 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_81
timestamp 1723858470
transform 1 0 552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1723858470
transform -1 0 23368 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_82
timestamp 1723858470
transform 1 0 552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1723858470
transform -1 0 23368 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_83
timestamp 1723858470
transform 1 0 552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1723858470
transform -1 0 23368 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1723858470
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1723858470
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1723858470
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1723858470
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_89
timestamp 1723858470
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_90
timestamp 1723858470
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_91
timestamp 1723858470
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1723858470
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1723858470
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_94
timestamp 1723858470
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_95
timestamp 1723858470
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1723858470
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1723858470
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1723858470
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1723858470
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1723858470
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1723858470
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1723858470
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1723858470
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_104
timestamp 1723858470
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1723858470
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1723858470
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1723858470
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_108
timestamp 1723858470
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_109
timestamp 1723858470
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_110
timestamp 1723858470
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1723858470
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_112
timestamp 1723858470
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_113
timestamp 1723858470
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_114
timestamp 1723858470
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_115
timestamp 1723858470
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1723858470
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_117
timestamp 1723858470
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_118
timestamp 1723858470
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_119
timestamp 1723858470
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1723858470
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1723858470
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1723858470
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_123
timestamp 1723858470
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1723858470
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1723858470
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1723858470
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1723858470
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1723858470
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1723858470
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1723858470
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1723858470
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp 1723858470
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp 1723858470
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1723858470
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1723858470
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_136
timestamp 1723858470
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_137
timestamp 1723858470
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_138
timestamp 1723858470
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1723858470
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_140
timestamp 1723858470
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_141
timestamp 1723858470
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_142
timestamp 1723858470
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_143
timestamp 1723858470
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_144
timestamp 1723858470
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_145
timestamp 1723858470
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_146
timestamp 1723858470
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_147
timestamp 1723858470
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_148
timestamp 1723858470
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_149
timestamp 1723858470
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_150
timestamp 1723858470
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_151
timestamp 1723858470
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_152
timestamp 1723858470
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_153
timestamp 1723858470
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_154
timestamp 1723858470
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_155
timestamp 1723858470
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp 1723858470
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_157
timestamp 1723858470
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_158
timestamp 1723858470
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_159
timestamp 1723858470
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp 1723858470
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp 1723858470
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_162
timestamp 1723858470
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_163
timestamp 1723858470
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp 1723858470
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp 1723858470
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_166
timestamp 1723858470
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_167
timestamp 1723858470
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp 1723858470
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp 1723858470
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_170
timestamp 1723858470
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_171
timestamp 1723858470
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp 1723858470
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp 1723858470
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_174
timestamp 1723858470
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_175
timestamp 1723858470
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_176
timestamp 1723858470
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp 1723858470
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_178
timestamp 1723858470
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_179
timestamp 1723858470
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_180
timestamp 1723858470
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_181
timestamp 1723858470
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_182
timestamp 1723858470
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_183
timestamp 1723858470
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_184
timestamp 1723858470
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_185
timestamp 1723858470
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_186
timestamp 1723858470
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_187
timestamp 1723858470
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_188
timestamp 1723858470
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_189
timestamp 1723858470
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_190
timestamp 1723858470
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_191
timestamp 1723858470
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_192
timestamp 1723858470
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_193
timestamp 1723858470
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_194
timestamp 1723858470
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_195
timestamp 1723858470
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_196
timestamp 1723858470
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_197
timestamp 1723858470
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_198
timestamp 1723858470
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_199
timestamp 1723858470
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_200
timestamp 1723858470
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_201
timestamp 1723858470
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_202
timestamp 1723858470
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_203
timestamp 1723858470
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_204
timestamp 1723858470
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_205
timestamp 1723858470
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_206
timestamp 1723858470
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_207
timestamp 1723858470
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_208
timestamp 1723858470
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_209
timestamp 1723858470
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_210
timestamp 1723858470
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_211
timestamp 1723858470
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_212
timestamp 1723858470
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_213
timestamp 1723858470
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_214
timestamp 1723858470
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_215
timestamp 1723858470
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_216
timestamp 1723858470
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_217
timestamp 1723858470
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_218
timestamp 1723858470
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_219
timestamp 1723858470
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_220
timestamp 1723858470
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_221
timestamp 1723858470
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_222
timestamp 1723858470
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_223
timestamp 1723858470
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_224
timestamp 1723858470
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_225
timestamp 1723858470
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_226
timestamp 1723858470
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_227
timestamp 1723858470
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_228
timestamp 1723858470
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_229
timestamp 1723858470
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_230
timestamp 1723858470
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_231
timestamp 1723858470
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_232
timestamp 1723858470
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_233
timestamp 1723858470
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_234
timestamp 1723858470
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_235
timestamp 1723858470
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_236
timestamp 1723858470
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_237
timestamp 1723858470
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_238
timestamp 1723858470
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_239
timestamp 1723858470
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_240
timestamp 1723858470
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_241
timestamp 1723858470
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_242
timestamp 1723858470
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_243
timestamp 1723858470
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_244
timestamp 1723858470
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_245
timestamp 1723858470
transform 1 0 10856 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_246
timestamp 1723858470
transform 1 0 16008 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_247
timestamp 1723858470
transform 1 0 21160 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_248
timestamp 1723858470
transform 1 0 3128 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_249
timestamp 1723858470
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_250
timestamp 1723858470
transform 1 0 13432 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_251
timestamp 1723858470
transform 1 0 18584 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_252
timestamp 1723858470
transform 1 0 3128 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_253
timestamp 1723858470
transform 1 0 5704 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_254
timestamp 1723858470
transform 1 0 8280 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_255
timestamp 1723858470
transform 1 0 10856 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_256
timestamp 1723858470
transform 1 0 13432 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_257
timestamp 1723858470
transform 1 0 16008 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_258
timestamp 1723858470
transform 1 0 18584 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_259
timestamp 1723858470
transform 1 0 21160 0 -1 23392
box -38 -48 130 592
<< labels >>
flabel metal4 s 4316 496 4636 23440 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3656 496 3976 23440 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 23600 3816 24000 3936 0 FreeSans 480 0 0 0 clk_in
port 2 nsew signal input
flabel metal3 s 23600 19592 24000 19712 0 FreeSans 480 0 0 0 clk_out
port 3 nsew signal output
flabel metal3 s 23600 11704 24000 11824 0 FreeSans 480 0 0 0 nrst
port 4 nsew signal input
flabel metal2 s 1674 23600 1730 24000 0 FreeSans 224 90 0 0 scale[0]
port 5 nsew signal input
flabel metal2 s 4618 23600 4674 24000 0 FreeSans 224 90 0 0 scale[1]
port 6 nsew signal input
flabel metal2 s 7562 23600 7618 24000 0 FreeSans 224 90 0 0 scale[2]
port 7 nsew signal input
flabel metal2 s 10506 23600 10562 24000 0 FreeSans 224 90 0 0 scale[3]
port 8 nsew signal input
flabel metal2 s 13450 23600 13506 24000 0 FreeSans 224 90 0 0 scale[4]
port 9 nsew signal input
flabel metal2 s 16394 23600 16450 24000 0 FreeSans 224 90 0 0 scale[5]
port 10 nsew signal input
flabel metal2 s 19338 23600 19394 24000 0 FreeSans 224 90 0 0 scale[6]
port 11 nsew signal input
flabel metal2 s 22282 23600 22338 24000 0 FreeSans 224 90 0 0 scale[7]
port 12 nsew signal input
rlabel metal1 11960 23392 11960 23392 0 VGND
rlabel metal1 11960 22848 11960 22848 0 VPWR
rlabel via1 6030 12750 6030 12750 0 _0000_
rlabel metal1 5872 15606 5872 15606 0 _0001_
rlabel metal1 5704 13498 5704 13498 0 _0002_
rlabel metal1 6956 13838 6956 13838 0 _0003_
rlabel metal1 7406 12954 7406 12954 0 _0004_
rlabel metal1 8965 12682 8965 12682 0 _0005_
rlabel metal2 9430 11458 9430 11458 0 _0006_
rlabel metal2 11270 11458 11270 11458 0 _0007_
rlabel via1 11633 12342 11633 12342 0 _0008_
rlabel metal1 12930 12750 12930 12750 0 _0009_
rlabel via1 14209 12750 14209 12750 0 _0010_
rlabel metal1 14250 12274 14250 12274 0 _0011_
rlabel metal1 15175 11662 15175 11662 0 _0012_
rlabel metal2 16146 13634 16146 13634 0 _0013_
rlabel metal1 16555 15606 16555 15606 0 _0014_
rlabel via1 16785 14926 16785 14926 0 _0015_
rlabel metal1 18896 17102 18896 17102 0 _0016_
rlabel metal1 18844 17782 18844 17782 0 _0017_
rlabel metal1 19913 18870 19913 18870 0 _0018_
rlabel metal2 21298 16898 21298 16898 0 _0019_
rlabel via1 22498 19278 22498 19278 0 _0020_
rlabel metal1 21420 18870 21420 18870 0 _0021_
rlabel metal1 5294 6902 5294 6902 0 _0022_
rlabel metal1 7007 6154 7007 6154 0 _0023_
rlabel metal1 6016 6834 6016 6834 0 _0024_
rlabel metal1 5366 7242 5366 7242 0 _0025_
rlabel metal1 5014 9690 5014 9690 0 _0026_
rlabel metal1 5096 9486 5096 9486 0 _0027_
rlabel metal2 6946 9894 6946 9894 0 _0028_
rlabel metal1 7488 9010 7488 9010 0 _0029_
rlabel via1 8974 7990 8974 7990 0 _0030_
rlabel metal2 9338 8194 9338 8194 0 _0031_
rlabel metal2 10442 7072 10442 7072 0 _0032_
rlabel metal1 11162 7990 11162 7990 0 _0033_
rlabel metal1 11628 8398 11628 8398 0 _0034_
rlabel metal1 13508 7990 13508 7990 0 _0035_
rlabel metal1 14020 8398 14020 8398 0 _0036_
rlabel metal2 15502 8194 15502 8194 0 _0037_
rlabel metal2 17618 8806 17618 8806 0 _0038_
rlabel metal2 17526 9860 17526 9860 0 _0039_
rlabel via1 18266 10574 18266 10574 0 _0040_
rlabel metal2 18262 12070 18262 12070 0 _0041_
rlabel via1 17981 12342 17981 12342 0 _0042_
rlabel metal1 19816 12750 19816 12750 0 _0043_
rlabel metal1 19810 11594 19810 11594 0 _0044_
rlabel metal2 21114 13396 21114 13396 0 _0045_
rlabel metal1 21834 12342 21834 12342 0 _0046_
rlabel metal2 21574 11458 21574 11458 0 _0047_
rlabel via1 21845 9486 21845 9486 0 _0048_
rlabel metal1 21466 9078 21466 9078 0 _0049_
rlabel metal1 21615 7990 21615 7990 0 _0050_
rlabel metal2 20194 9282 20194 9282 0 _0051_
rlabel via1 19177 8398 19177 8398 0 _0052_
rlabel metal1 18804 9010 18804 9010 0 _0053_
rlabel metal1 21840 18190 21840 18190 0 _0054_
rlabel metal2 21942 18258 21942 18258 0 _0055_
rlabel metal1 21390 18394 21390 18394 0 _0056_
rlabel metal1 5750 17136 5750 17136 0 _0057_
rlabel metal1 5566 17714 5566 17714 0 _0058_
rlabel metal1 8694 21522 8694 21522 0 _0059_
rlabel metal1 16468 21454 16468 21454 0 _0060_
rlabel metal2 7130 12444 7130 12444 0 _0061_
rlabel via1 7498 11730 7498 11730 0 _0062_
rlabel metal2 9522 10880 9522 10880 0 _0063_
rlabel metal2 12558 10982 12558 10982 0 _0064_
rlabel metal1 11224 10574 11224 10574 0 _0065_
rlabel metal2 15318 11356 15318 11356 0 _0066_
rlabel metal2 14582 10812 14582 10812 0 _0067_
rlabel metal1 16882 13838 16882 13838 0 _0068_
rlabel metal1 17940 14858 17940 14858 0 _0069_
rlabel metal1 19366 16082 19366 16082 0 _0070_
rlabel metal2 19734 15708 19734 15708 0 _0071_
rlabel metal1 20332 15334 20332 15334 0 _0072_
rlabel metal1 22356 14518 22356 14518 0 _0073_
rlabel metal1 22954 14348 22954 14348 0 _0074_
rlabel metal1 5014 16762 5014 16762 0 _0075_
rlabel metal2 5106 15844 5106 15844 0 _0076_
rlabel metal1 5336 21318 5336 21318 0 _0077_
rlabel metal2 5106 20672 5106 20672 0 _0078_
rlabel via1 5474 20570 5474 20570 0 _0079_
rlabel metal1 5566 20298 5566 20298 0 _0080_
rlabel metal1 5566 17782 5566 17782 0 _0081_
rlabel metal1 9062 21488 9062 21488 0 _0082_
rlabel metal2 7682 16983 7682 16983 0 _0083_
rlabel metal1 10074 21556 10074 21556 0 _0084_
rlabel metal2 9706 21454 9706 21454 0 _0085_
rlabel metal1 9292 21386 9292 21386 0 _0086_
rlabel metal1 8234 12682 8234 12682 0 _0087_
rlabel metal1 12466 22032 12466 22032 0 _0088_
rlabel metal1 9890 20978 9890 20978 0 _0089_
rlabel metal1 7728 22950 7728 22950 0 _0090_
rlabel metal2 11178 21420 11178 21420 0 _0091_
rlabel metal1 9246 14926 9246 14926 0 _0092_
rlabel metal1 11086 22134 11086 22134 0 _0093_
rlabel metal1 9108 19890 9108 19890 0 _0094_
rlabel metal1 8188 20366 8188 20366 0 _0095_
rlabel metal2 7498 17748 7498 17748 0 _0096_
rlabel metal1 6256 17714 6256 17714 0 _0097_
rlabel metal1 7314 18836 7314 18836 0 _0098_
rlabel metal2 8786 18564 8786 18564 0 _0099_
rlabel metal2 8326 19380 8326 19380 0 _0100_
rlabel metal2 9890 17374 9890 17374 0 _0101_
rlabel metal2 9522 19244 9522 19244 0 _0102_
rlabel via1 10074 17510 10074 17510 0 _0103_
rlabel via1 9430 14926 9430 14926 0 _0104_
rlabel metal2 9798 14314 9798 14314 0 _0105_
rlabel metal2 9246 14722 9246 14722 0 _0106_
rlabel metal1 9522 14450 9522 14450 0 _0107_
rlabel metal1 9844 14314 9844 14314 0 _0108_
rlabel metal1 10028 13294 10028 13294 0 _0109_
rlabel metal2 9614 13702 9614 13702 0 _0110_
rlabel metal2 12006 20400 12006 20400 0 _0111_
rlabel metal2 10810 15844 10810 15844 0 _0112_
rlabel metal1 9798 19244 9798 19244 0 _0113_
rlabel metal1 10856 18394 10856 18394 0 _0114_
rlabel metal1 6210 18156 6210 18156 0 _0115_
rlabel metal1 6716 17714 6716 17714 0 _0116_
rlabel metal1 6486 17646 6486 17646 0 _0117_
rlabel metal1 9246 17102 9246 17102 0 _0118_
rlabel metal1 8602 17748 8602 17748 0 _0119_
rlabel metal1 9982 17000 9982 17000 0 _0120_
rlabel metal2 9706 14705 9706 14705 0 _0121_
rlabel metal2 10258 15436 10258 15436 0 _0122_
rlabel metal2 9982 14042 9982 14042 0 _0123_
rlabel metal1 9982 13396 9982 13396 0 _0124_
rlabel metal1 8786 13430 8786 13430 0 _0125_
rlabel via1 9338 13226 9338 13226 0 _0126_
rlabel metal2 9890 11696 9890 11696 0 _0127_
rlabel metal1 10120 17646 10120 17646 0 _0128_
rlabel metal1 7866 19924 7866 19924 0 _0129_
rlabel metal2 5474 16898 5474 16898 0 _0130_
rlabel metal1 6946 16490 6946 16490 0 _0131_
rlabel metal2 7314 18700 7314 18700 0 _0132_
rlabel metal2 7130 16422 7130 16422 0 _0133_
rlabel metal2 7774 16014 7774 16014 0 _0134_
rlabel metal1 7682 16150 7682 16150 0 _0135_
rlabel metal1 9522 16082 9522 16082 0 _0136_
rlabel metal1 9246 16082 9246 16082 0 _0137_
rlabel metal2 11914 15470 11914 15470 0 _0138_
rlabel metal1 10903 15980 10903 15980 0 _0139_
rlabel metal2 12006 15708 12006 15708 0 _0140_
rlabel metal1 10028 14450 10028 14450 0 _0141_
rlabel metal2 11362 14688 11362 14688 0 _0142_
rlabel metal2 10626 14314 10626 14314 0 _0143_
rlabel metal2 10442 13226 10442 13226 0 _0144_
rlabel metal1 10258 12818 10258 12818 0 _0145_
rlabel metal1 11270 12614 11270 12614 0 _0146_
rlabel metal1 16698 19890 16698 19890 0 _0147_
rlabel metal1 5796 20978 5796 20978 0 _0148_
rlabel metal1 12006 22202 12006 22202 0 _0149_
rlabel metal2 6394 17170 6394 17170 0 _0150_
rlabel metal2 6118 16762 6118 16762 0 _0151_
rlabel metal2 6946 16694 6946 16694 0 _0152_
rlabel metal1 7314 16082 7314 16082 0 _0153_
rlabel metal2 8142 15708 8142 15708 0 _0154_
rlabel metal1 8050 15436 8050 15436 0 _0155_
rlabel metal1 12696 15538 12696 15538 0 _0156_
rlabel metal1 10948 15470 10948 15470 0 _0157_
rlabel metal2 12558 15334 12558 15334 0 _0158_
rlabel metal1 11914 14926 11914 14926 0 _0159_
rlabel metal1 13662 14824 13662 14824 0 _0160_
rlabel metal2 11638 14892 11638 14892 0 _0161_
rlabel metal2 13202 14246 13202 14246 0 _0162_
rlabel metal1 11270 14552 11270 14552 0 _0163_
rlabel metal1 10864 14790 10864 14790 0 _0164_
rlabel metal1 11592 14382 11592 14382 0 _0165_
rlabel metal1 12834 14416 12834 14416 0 _0166_
rlabel metal2 11822 13804 11822 13804 0 _0167_
rlabel metal1 12006 12954 12006 12954 0 _0168_
rlabel metal1 17066 22066 17066 22066 0 _0169_
rlabel metal2 16146 21726 16146 21726 0 _0170_
rlabel metal1 16606 21556 16606 21556 0 _0171_
rlabel metal1 13340 22066 13340 22066 0 _0172_
rlabel metal1 17296 21658 17296 21658 0 _0173_
rlabel metal1 16514 20944 16514 20944 0 _0174_
rlabel metal2 11776 22066 11776 22066 0 _0175_
rlabel metal1 12006 22576 12006 22576 0 _0176_
rlabel metal1 12788 22202 12788 22202 0 _0177_
rlabel metal1 12374 22542 12374 22542 0 _0178_
rlabel metal2 13110 21828 13110 21828 0 _0179_
rlabel metal2 13018 18938 13018 18938 0 _0180_
rlabel metal1 13202 16116 13202 16116 0 _0181_
rlabel metal1 13616 15946 13616 15946 0 _0182_
rlabel metal1 12880 16082 12880 16082 0 _0183_
rlabel metal1 12880 15538 12880 15538 0 _0184_
rlabel metal2 13570 15130 13570 15130 0 _0185_
rlabel metal1 13478 15062 13478 15062 0 _0186_
rlabel metal1 13938 14450 13938 14450 0 _0187_
rlabel metal2 13754 13600 13754 13600 0 _0188_
rlabel metal2 12834 13532 12834 13532 0 _0189_
rlabel metal1 14674 13294 14674 13294 0 _0190_
rlabel metal2 18906 21386 18906 21386 0 _0191_
rlabel metal1 20194 23222 20194 23222 0 _0192_
rlabel metal1 19136 22066 19136 22066 0 _0193_
rlabel metal2 20010 22780 20010 22780 0 _0194_
rlabel metal1 18722 21998 18722 21998 0 _0195_
rlabel metal1 13202 21488 13202 21488 0 _0196_
rlabel metal1 13110 21522 13110 21522 0 _0197_
rlabel metal1 13386 22610 13386 22610 0 _0198_
rlabel metal1 13570 21590 13570 21590 0 _0199_
rlabel metal1 13478 20978 13478 20978 0 _0200_
rlabel metal2 14122 21216 14122 21216 0 _0201_
rlabel metal1 14260 21454 14260 21454 0 _0202_
rlabel metal2 14674 21046 14674 21046 0 _0203_
rlabel metal1 15226 15946 15226 15946 0 _0204_
rlabel metal1 14950 16082 14950 16082 0 _0205_
rlabel metal1 15088 16218 15088 16218 0 _0206_
rlabel metal1 13892 15130 13892 15130 0 _0207_
rlabel metal2 14306 13804 14306 13804 0 _0208_
rlabel metal1 14214 13362 14214 13362 0 _0209_
rlabel metal1 15226 16558 15226 16558 0 _0210_
rlabel metal1 21390 21386 21390 21386 0 _0211_
rlabel metal1 13570 20502 13570 20502 0 _0212_
rlabel metal1 10534 20978 10534 20978 0 _0213_
rlabel metal1 10672 21318 10672 21318 0 _0214_
rlabel metal2 9246 21760 9246 21760 0 _0215_
rlabel metal1 10718 21488 10718 21488 0 _0216_
rlabel metal1 10442 21420 10442 21420 0 _0217_
rlabel metal2 14122 22015 14122 22015 0 _0218_
rlabel metal1 14582 22576 14582 22576 0 _0219_
rlabel metal1 15226 22202 15226 22202 0 _0220_
rlabel metal2 15042 21488 15042 21488 0 _0221_
rlabel metal2 15042 16915 15042 16915 0 _0222_
rlabel metal2 15502 16456 15502 16456 0 _0223_
rlabel metal1 14674 16592 14674 16592 0 _0224_
rlabel metal2 14398 15402 14398 15402 0 _0225_
rlabel metal1 14490 13838 14490 13838 0 _0226_
rlabel metal2 14674 14144 14674 14144 0 _0227_
rlabel metal1 13800 12274 13800 12274 0 _0228_
rlabel metal2 8970 19516 8970 19516 0 _0229_
rlabel metal1 10212 18938 10212 18938 0 _0230_
rlabel metal2 12466 20128 12466 20128 0 _0231_
rlabel metal1 12834 20400 12834 20400 0 _0232_
rlabel metal2 13662 20094 13662 20094 0 _0233_
rlabel metal1 13524 19822 13524 19822 0 _0234_
rlabel metal2 13846 20060 13846 20060 0 _0235_
rlabel metal1 14214 19958 14214 19958 0 _0236_
rlabel metal1 14582 19822 14582 19822 0 _0237_
rlabel metal1 14904 18938 14904 18938 0 _0238_
rlabel metal1 14858 19686 14858 19686 0 _0239_
rlabel metal2 14674 16116 14674 16116 0 _0240_
rlabel metal1 15088 17102 15088 17102 0 _0241_
rlabel metal1 14950 18258 14950 18258 0 _0242_
rlabel metal1 15732 12818 15732 12818 0 _0243_
rlabel metal1 10672 18190 10672 18190 0 _0244_
rlabel metal1 10902 18292 10902 18292 0 _0245_
rlabel metal2 11638 18394 11638 18394 0 _0246_
rlabel metal2 12006 18462 12006 18462 0 _0247_
rlabel metal1 13938 18700 13938 18700 0 _0248_
rlabel metal2 14582 18836 14582 18836 0 _0249_
rlabel metal1 14076 18802 14076 18802 0 _0250_
rlabel metal1 14352 19754 14352 19754 0 _0251_
rlabel metal2 14766 18972 14766 18972 0 _0252_
rlabel metal1 14536 18734 14536 18734 0 _0253_
rlabel metal1 16514 13294 16514 13294 0 _0254_
rlabel metal1 5474 18734 5474 18734 0 _0255_
rlabel metal2 6762 18428 6762 18428 0 _0256_
rlabel metal1 7406 18394 7406 18394 0 _0257_
rlabel metal2 7222 17952 7222 17952 0 _0258_
rlabel metal1 11178 17748 11178 17748 0 _0259_
rlabel metal1 10626 17170 10626 17170 0 _0260_
rlabel metal1 11408 17646 11408 17646 0 _0261_
rlabel metal2 12374 17476 12374 17476 0 _0262_
rlabel metal1 13386 17748 13386 17748 0 _0263_
rlabel metal2 13294 17986 13294 17986 0 _0264_
rlabel metal1 16514 16966 16514 16966 0 _0265_
rlabel metal2 17434 17510 17434 17510 0 _0266_
rlabel metal1 16008 17782 16008 17782 0 _0267_
rlabel metal2 15594 17612 15594 17612 0 _0268_
rlabel metal1 15548 16626 15548 16626 0 _0269_
rlabel metal1 16330 17544 16330 17544 0 _0270_
rlabel metal1 17066 16660 17066 16660 0 _0271_
rlabel metal2 16146 16218 16146 16218 0 _0272_
rlabel metal2 16330 20740 16330 20740 0 _0273_
rlabel metal2 6670 20570 6670 20570 0 _0274_
rlabel metal1 6808 19890 6808 19890 0 _0275_
rlabel metal1 6578 19788 6578 19788 0 _0276_
rlabel metal1 7406 19482 7406 19482 0 _0277_
rlabel metal1 7406 19754 7406 19754 0 _0278_
rlabel metal1 15410 19380 15410 19380 0 _0279_
rlabel metal2 15502 19023 15502 19023 0 _0280_
rlabel metal1 16422 19210 16422 19210 0 _0281_
rlabel metal2 16330 19006 16330 19006 0 _0282_
rlabel metal1 16008 18190 16008 18190 0 _0283_
rlabel metal1 15778 17680 15778 17680 0 _0284_
rlabel metal1 16376 17714 16376 17714 0 _0285_
rlabel metal1 16974 17714 16974 17714 0 _0286_
rlabel metal1 16928 17102 16928 17102 0 _0287_
rlabel metal2 17158 17544 17158 17544 0 _0288_
rlabel metal2 16974 16626 16974 16626 0 _0289_
rlabel metal2 17066 16218 17066 16218 0 _0290_
rlabel metal2 16514 21556 16514 21556 0 _0291_
rlabel metal1 18078 21488 18078 21488 0 _0292_
rlabel metal2 17618 21488 17618 21488 0 _0293_
rlabel metal1 17940 21454 17940 21454 0 _0294_
rlabel metal2 17342 21284 17342 21284 0 _0295_
rlabel metal1 17434 20366 17434 20366 0 _0296_
rlabel metal1 17250 20366 17250 20366 0 _0297_
rlabel metal2 18170 20128 18170 20128 0 _0298_
rlabel metal2 17158 20060 17158 20060 0 _0299_
rlabel metal1 18078 19924 18078 19924 0 _0300_
rlabel metal2 17986 19516 17986 19516 0 _0301_
rlabel metal1 18078 19244 18078 19244 0 _0302_
rlabel via1 18722 19482 18722 19482 0 _0303_
rlabel metal1 18814 18836 18814 18836 0 _0304_
rlabel metal1 18676 18190 18676 18190 0 _0305_
rlabel metal1 14766 15062 14766 15062 0 _0306_
rlabel metal1 15778 17238 15778 17238 0 _0307_
rlabel metal1 17296 17170 17296 17170 0 _0308_
rlabel metal2 17710 17748 17710 17748 0 _0309_
rlabel metal2 17618 17612 17618 17612 0 _0310_
rlabel metal1 18170 17102 18170 17102 0 _0311_
rlabel metal1 18860 18258 18860 18258 0 _0312_
rlabel metal1 18400 16490 18400 16490 0 _0313_
rlabel metal1 18676 16762 18676 16762 0 _0314_
rlabel metal1 18308 22202 18308 22202 0 _0315_
rlabel metal1 19540 21386 19540 21386 0 _0316_
rlabel metal2 18814 22338 18814 22338 0 _0317_
rlabel metal1 19044 21522 19044 21522 0 _0318_
rlabel metal1 19366 21420 19366 21420 0 _0319_
rlabel via1 19266 20026 19266 20026 0 _0320_
rlabel metal1 18998 19278 18998 19278 0 _0321_
rlabel metal2 18354 20060 18354 20060 0 _0322_
rlabel metal1 18492 18734 18492 18734 0 _0323_
rlabel metal2 18538 18190 18538 18190 0 _0324_
rlabel metal2 18722 17884 18722 17884 0 _0325_
rlabel metal1 21758 22746 21758 22746 0 _0326_
rlabel metal2 22586 22542 22586 22542 0 _0327_
rlabel metal1 22310 22134 22310 22134 0 _0328_
rlabel metal1 22172 22474 22172 22474 0 _0329_
rlabel metal1 22218 21896 22218 21896 0 _0330_
rlabel metal1 22034 21488 22034 21488 0 _0331_
rlabel metal1 20746 21488 20746 21488 0 _0332_
rlabel metal1 20117 21454 20117 21454 0 _0333_
rlabel metal1 21298 20978 21298 20978 0 _0334_
rlabel metal2 20470 21148 20470 21148 0 _0335_
rlabel metal2 20286 20332 20286 20332 0 _0336_
rlabel metal2 19826 19142 19826 19142 0 _0337_
rlabel metal2 18538 20060 18538 20060 0 _0338_
rlabel metal1 19734 19856 19734 19856 0 _0339_
rlabel metal1 21436 20570 21436 20570 0 _0340_
rlabel metal1 20240 19346 20240 19346 0 _0341_
rlabel metal1 20424 18394 20424 18394 0 _0342_
rlabel metal2 21758 19516 21758 19516 0 _0343_
rlabel metal1 21390 22134 21390 22134 0 _0344_
rlabel metal2 21758 21420 21758 21420 0 _0345_
rlabel metal2 22126 21352 22126 21352 0 _0346_
rlabel metal1 21482 20366 21482 20366 0 _0347_
rlabel metal2 22678 20094 22678 20094 0 _0348_
rlabel metal1 22586 19890 22586 19890 0 _0349_
rlabel metal2 22770 18190 22770 18190 0 _0350_
rlabel metal2 21298 20400 21298 20400 0 _0351_
rlabel metal1 22080 19958 22080 19958 0 _0352_
rlabel metal1 21574 19890 21574 19890 0 _0353_
rlabel metal1 22310 8602 22310 8602 0 _0354_
rlabel metal2 22770 12614 22770 12614 0 _0355_
rlabel metal1 22448 14450 22448 14450 0 _0356_
rlabel metal1 22172 14450 22172 14450 0 _0357_
rlabel metal1 21022 10030 21022 10030 0 _0358_
rlabel metal1 21390 10234 21390 10234 0 _0359_
rlabel metal2 21942 14212 21942 14212 0 _0360_
rlabel metal2 22402 15130 22402 15130 0 _0361_
rlabel metal2 21298 15164 21298 15164 0 _0362_
rlabel metal1 21988 15062 21988 15062 0 _0363_
rlabel metal1 20391 15674 20391 15674 0 _0364_
rlabel metal1 20792 15538 20792 15538 0 _0365_
rlabel metal2 20654 15232 20654 15232 0 _0366_
rlabel metal2 19918 15708 19918 15708 0 _0367_
rlabel metal2 19826 15164 19826 15164 0 _0368_
rlabel metal1 20516 14994 20516 14994 0 _0369_
rlabel metal2 18446 14858 18446 14858 0 _0370_
rlabel metal1 19044 13838 19044 13838 0 _0371_
rlabel metal2 17756 14450 17756 14450 0 _0372_
rlabel metal1 18998 14586 18998 14586 0 _0373_
rlabel metal1 18127 14586 18127 14586 0 _0374_
rlabel metal2 19090 14416 19090 14416 0 _0375_
rlabel metal2 18354 14076 18354 14076 0 _0376_
rlabel metal2 17986 14246 17986 14246 0 _0377_
rlabel metal1 17802 14416 17802 14416 0 _0378_
rlabel metal1 18538 13906 18538 13906 0 _0379_
rlabel metal2 16882 11594 16882 11594 0 _0380_
rlabel metal2 17434 11492 17434 11492 0 _0381_
rlabel metal1 15686 11254 15686 11254 0 _0382_
rlabel metal2 16790 11594 16790 11594 0 _0383_
rlabel metal1 16606 11050 16606 11050 0 _0384_
rlabel metal2 15134 10234 15134 10234 0 _0385_
rlabel metal2 15318 9690 15318 9690 0 _0386_
rlabel metal1 15042 10574 15042 10574 0 _0387_
rlabel metal1 14720 10030 14720 10030 0 _0388_
rlabel metal2 14858 9792 14858 9792 0 _0389_
rlabel metal1 13570 10540 13570 10540 0 _0390_
rlabel metal2 13754 10234 13754 10234 0 _0391_
rlabel metal1 14720 9962 14720 9962 0 _0392_
rlabel metal2 12190 9996 12190 9996 0 _0393_
rlabel metal2 12466 9860 12466 9860 0 _0394_
rlabel metal2 11546 10778 11546 10778 0 _0395_
rlabel metal2 11638 10234 11638 10234 0 _0396_
rlabel metal1 12098 9894 12098 9894 0 _0397_
rlabel metal1 10626 9554 10626 9554 0 _0398_
rlabel metal1 11822 9690 11822 9690 0 _0399_
rlabel metal1 9392 10438 9392 10438 0 _0400_
rlabel metal2 9706 10268 9706 10268 0 _0401_
rlabel metal1 10074 9894 10074 9894 0 _0402_
rlabel metal2 8878 10336 8878 10336 0 _0403_
rlabel metal1 9154 9996 9154 9996 0 _0404_
rlabel metal2 7406 11628 7406 11628 0 _0405_
rlabel metal1 7866 11084 7866 11084 0 _0406_
rlabel metal1 7728 10982 7728 10982 0 _0407_
rlabel metal2 7222 12036 7222 12036 0 _0408_
rlabel metal2 6854 11356 6854 11356 0 _0409_
rlabel metal1 6900 10982 6900 10982 0 _0410_
rlabel metal2 5842 11900 5842 11900 0 _0411_
rlabel metal1 6624 11186 6624 11186 0 _0412_
rlabel metal1 7636 6970 7636 6970 0 _0413_
rlabel metal2 4462 7752 4462 7752 0 _0414_
rlabel metal1 5014 7378 5014 7378 0 _0415_
rlabel metal1 5152 10982 5152 10982 0 _0416_
rlabel metal1 6315 11322 6315 11322 0 _0417_
rlabel metal1 6440 11254 6440 11254 0 _0418_
rlabel metal1 7774 11152 7774 11152 0 _0419_
rlabel metal1 9384 10166 9384 10166 0 _0420_
rlabel metal1 12190 10200 12190 10200 0 _0421_
rlabel metal1 14904 9486 14904 9486 0 _0422_
rlabel metal1 16054 9622 16054 9622 0 _0423_
rlabel metal1 18170 11798 18170 11798 0 _0424_
rlabel metal1 19918 14042 19918 14042 0 _0425_
rlabel metal2 22034 15164 22034 15164 0 _0426_
rlabel metal1 22218 14994 22218 14994 0 _0427_
rlabel metal2 22494 14552 22494 14552 0 _0428_
rlabel metal1 22241 13362 22241 13362 0 _0429_
rlabel metal1 22724 13362 22724 13362 0 _0430_
rlabel metal1 7528 7242 7528 7242 0 _0431_
rlabel metal1 5720 7990 5720 7990 0 _0432_
rlabel metal1 5060 7242 5060 7242 0 _0433_
rlabel metal1 4692 9690 4692 9690 0 _0434_
rlabel metal2 5290 9282 5290 9282 0 _0435_
rlabel metal1 5382 10234 5382 10234 0 _0436_
rlabel metal1 4830 9928 4830 9928 0 _0437_
rlabel metal1 6026 9486 6026 9486 0 _0438_
rlabel metal2 6762 10064 6762 10064 0 _0439_
rlabel metal2 7130 8704 7130 8704 0 _0440_
rlabel metal1 7373 9146 7373 9146 0 _0441_
rlabel metal2 8418 9044 8418 9044 0 _0442_
rlabel metal2 9982 9418 9982 9418 0 _0443_
rlabel metal1 11492 9146 11492 9146 0 _0444_
rlabel metal2 9522 8534 9522 8534 0 _0445_
rlabel metal1 10442 6630 10442 6630 0 _0446_
rlabel via1 10618 6970 10618 6970 0 _0447_
rlabel metal1 10994 8908 10994 8908 0 _0448_
rlabel metal2 10350 8330 10350 8330 0 _0449_
rlabel metal2 14950 8160 14950 8160 0 _0450_
rlabel metal2 12466 8704 12466 8704 0 _0451_
rlabel metal1 13432 8602 13432 8602 0 _0452_
rlabel metal1 13356 8330 13356 8330 0 _0453_
rlabel metal2 14490 9316 14490 9316 0 _0454_
rlabel metal2 14122 8160 14122 8160 0 _0455_
rlabel metal1 17840 9418 17840 9418 0 _0456_
rlabel metal2 15318 8262 15318 8262 0 _0457_
rlabel metal1 17158 8602 17158 8602 0 _0458_
rlabel metal1 17396 8330 17396 8330 0 _0459_
rlabel metal1 16836 9622 16836 9622 0 _0460_
rlabel metal1 17066 9690 17066 9690 0 _0461_
rlabel metal1 17710 12784 17710 12784 0 _0462_
rlabel metal1 17710 10778 17710 10778 0 _0463_
rlabel metal1 17940 12682 17940 12682 0 _0464_
rlabel metal1 18040 11594 18040 11594 0 _0465_
rlabel metal1 20792 13294 20792 13294 0 _0466_
rlabel metal1 18446 12954 18446 12954 0 _0467_
rlabel metal1 20838 13362 20838 13362 0 _0468_
rlabel metal2 19918 13430 19918 13430 0 _0469_
rlabel metal1 20470 11322 20470 11322 0 _0470_
rlabel metal1 19780 11322 19780 11322 0 _0471_
rlabel metal1 22241 12682 22241 12682 0 _0472_
rlabel metal2 21298 13056 21298 13056 0 _0473_
rlabel metal2 22310 12308 22310 12308 0 _0474_
rlabel metal1 22356 12954 22356 12954 0 _0475_
rlabel metal2 22126 12172 22126 12172 0 _0476_
rlabel metal1 21988 10982 21988 10982 0 _0477_
rlabel metal2 22494 10268 22494 10268 0 _0478_
rlabel metal1 22540 9894 22540 9894 0 _0479_
rlabel metal1 21482 10540 21482 10540 0 _0480_
rlabel metal1 21896 10574 21896 10574 0 _0481_
rlabel metal2 21206 7956 21206 7956 0 _0482_
rlabel metal2 20470 8840 20470 8840 0 _0483_
rlabel metal1 20516 9010 20516 9010 0 _0484_
rlabel metal2 19734 8704 19734 8704 0 _0485_
rlabel metal2 19642 8738 19642 8738 0 _0486_
rlabel metal1 18860 8058 18860 8058 0 _0487_
rlabel metal1 18643 9146 18643 9146 0 _0488_
rlabel metal1 21620 17850 21620 17850 0 _0489_
rlabel metal2 23046 3961 23046 3961 0 clk_in
rlabel metal2 23046 18717 23046 18717 0 clk_out
rlabel metal2 4278 7140 4278 7140 0 count\[0\]
rlabel metal1 10810 7990 10810 7990 0 count\[10\]
rlabel metal2 11638 8534 11638 8534 0 count\[11\]
rlabel metal2 12834 8806 12834 8806 0 count\[12\]
rlabel metal1 14030 9418 14030 9418 0 count\[13\]
rlabel via1 14766 8262 14766 8262 0 count\[14\]
rlabel metal2 15410 9588 15410 9588 0 count\[15\]
rlabel metal1 16192 11254 16192 11254 0 count\[16\]
rlabel metal1 17388 11186 17388 11186 0 count\[17\]
rlabel metal1 17848 13838 17848 13838 0 count\[18\]
rlabel via1 17894 13430 17894 13430 0 count\[19\]
rlabel metal1 4554 7242 4554 7242 0 count\[1\]
rlabel metal1 18584 13158 18584 13158 0 count\[20\]
rlabel metal1 20010 13838 20010 13838 0 count\[21\]
rlabel metal1 20838 14858 20838 14858 0 count\[22\]
rlabel metal1 21620 14042 21620 14042 0 count\[23\]
rlabel metal1 23000 12070 23000 12070 0 count\[24\]
rlabel metal2 22402 11356 22402 11356 0 count\[25\]
rlabel metal1 22816 9350 22816 9350 0 count\[26\]
rlabel metal1 22402 10744 22402 10744 0 count\[27\]
rlabel metal1 20884 8262 20884 8262 0 count\[28\]
rlabel metal1 21022 9690 21022 9690 0 count\[29\]
rlabel metal1 5290 7922 5290 7922 0 count\[2\]
rlabel metal1 20608 10098 20608 10098 0 count\[30\]
rlabel metal1 21666 8330 21666 8330 0 count\[31\]
rlabel metal1 6486 7514 6486 7514 0 count\[3\]
rlabel metal1 5290 9078 5290 9078 0 count\[4\]
rlabel metal1 5014 10098 5014 10098 0 count\[5\]
rlabel metal1 6486 11628 6486 11628 0 count\[6\]
rlabel metal2 8602 11390 8602 11390 0 count\[7\]
rlabel metal1 7958 8602 7958 8602 0 count\[8\]
rlabel metal1 9338 10540 9338 10540 0 count\[9\]
rlabel metal1 18354 9112 18354 9112 0 net1
rlabel metal1 22586 23052 22586 23052 0 net10
rlabel metal1 9752 7990 9752 7990 0 net11
rlabel metal1 20700 8806 20700 8806 0 net12
rlabel metal1 20378 12682 20378 12682 0 net13
rlabel metal2 22678 12750 22678 12750 0 net14
rlabel metal1 20424 19346 20424 19346 0 net15
rlabel metal1 20608 19278 20608 19278 0 net16
rlabel metal2 12742 21726 12742 21726 0 net17
rlabel metal2 5290 18207 5290 18207 0 net18
rlabel metal2 5290 21726 5290 21726 0 net19
rlabel metal1 22448 17102 22448 17102 0 net2
rlabel via1 5566 16014 5566 16014 0 net20
rlabel metal2 22402 19414 22402 19414 0 net21
rlabel metal1 22310 17306 22310 17306 0 net22
rlabel metal1 8648 12750 8648 12750 0 net23
rlabel metal1 13340 7854 13340 7854 0 net24
rlabel metal2 13110 8500 13110 8500 0 net25
rlabel metal2 19228 12580 19228 12580 0 net26
rlabel metal1 21574 11662 21574 11662 0 net27
rlabel metal1 22586 17646 22586 17646 0 net28
rlabel metal1 20194 13906 20194 13906 0 net29
rlabel metal1 1978 23256 1978 23256 0 net3
rlabel metal1 5704 22066 5704 22066 0 net4
rlabel metal1 6900 20978 6900 20978 0 net5
rlabel metal1 6394 21488 6394 21488 0 net6
rlabel metal1 21758 23120 21758 23120 0 net7
rlabel metal2 17526 22712 17526 22712 0 net8
rlabel metal1 12834 19244 12834 19244 0 net9
rlabel metal2 23046 12257 23046 12257 0 nrst
rlabel metal2 1794 23443 1794 23443 0 scale[0]
rlabel metal2 4738 23443 4738 23443 0 scale[1]
rlabel metal1 8050 23188 8050 23188 0 scale[2]
rlabel metal2 10442 23477 10442 23477 0 scale[3]
rlabel metal2 13570 23443 13570 23443 0 scale[4]
rlabel metal1 16468 23154 16468 23154 0 scale[5]
rlabel metal2 19550 23477 19550 23477 0 scale[6]
rlabel metal1 22356 23154 22356 23154 0 scale[7]
rlabel metal1 22724 18054 22724 18054 0 signal_clk_out
rlabel metal1 9476 12614 9476 12614 0 true_scale\[10\]
rlabel metal2 10350 11322 10350 11322 0 true_scale\[11\]
rlabel metal1 12650 11118 12650 11118 0 true_scale\[12\]
rlabel metal1 12696 12410 12696 12410 0 true_scale\[13\]
rlabel metal2 12558 12954 12558 12954 0 true_scale\[14\]
rlabel metal2 15318 13124 15318 13124 0 true_scale\[15\]
rlabel metal1 14766 12070 14766 12070 0 true_scale\[16\]
rlabel metal1 15916 11866 15916 11866 0 true_scale\[17\]
rlabel metal1 16560 13430 16560 13430 0 true_scale\[18\]
rlabel metal2 17526 15810 17526 15810 0 true_scale\[19\]
rlabel metal2 17710 15776 17710 15776 0 true_scale\[20\]
rlabel metal2 20102 16490 20102 16490 0 true_scale\[21\]
rlabel metal1 19320 17510 19320 17510 0 true_scale\[22\]
rlabel metal1 20838 18258 20838 18258 0 true_scale\[23\]
rlabel metal2 21758 16796 21758 16796 0 true_scale\[24\]
rlabel metal2 22310 18054 22310 18054 0 true_scale\[25\]
rlabel metal1 22632 18938 22632 18938 0 true_scale\[26\]
rlabel metal1 5244 12614 5244 12614 0 true_scale\[5\]
rlabel metal1 6302 15334 6302 15334 0 true_scale\[6\]
rlabel metal2 6210 13770 6210 13770 0 true_scale\[7\]
rlabel metal1 7176 13770 7176 13770 0 true_scale\[8\]
rlabel metal1 8142 12750 8142 12750 0 true_scale\[9\]
<< properties >>
string FIXED_BBOX 0 0 24000 24000
<< end >>
