magic
tech sky130A
magscale 1 2
timestamp 1729368920
<< psubdiff >>
rect 2271 17263 2331 17297
rect 29791 17263 29851 17297
rect 2271 17237 2305 17263
rect 2271 1727 2305 1753
rect 29817 17237 29851 17263
rect 29817 1727 29851 1753
rect 2271 1693 2331 1727
rect 29791 1693 29851 1727
<< psubdiffcont >>
rect 2331 17263 29791 17297
rect 2271 1753 2305 17237
rect 29817 1753 29851 17237
rect 2331 1693 29791 1727
<< locali >>
rect 2271 17263 2331 17297
rect 29791 17263 29851 17297
rect 2271 17237 2305 17263
rect 2271 1727 2305 1753
rect 29817 17237 29851 17263
rect 29817 1727 29851 1753
rect 2271 1693 2331 1727
rect 29791 1693 29851 1727
<< metal1 >>
rect 5910 44690 5966 44720
rect 5896 44626 5906 44690
rect 5972 44682 5982 44690
rect 27650 44682 27660 44684
rect 5972 44626 27660 44682
rect 27724 44626 27734 44684
rect 8854 44538 8910 44570
rect 8836 44466 8846 44538
rect 8920 44532 8930 44538
rect 27116 44532 27126 44534
rect 8920 44476 27126 44532
rect 27190 44476 27200 44534
rect 8920 44466 8930 44476
rect 11798 44380 26628 44382
rect 11784 44308 11794 44380
rect 11868 44376 26628 44380
rect 11868 44326 26558 44376
rect 11868 44308 11878 44326
rect 26536 44318 26558 44326
rect 26622 44318 26632 44376
rect 11798 44302 11854 44308
rect 14742 44228 14798 44230
rect 14742 44214 14800 44228
rect 14734 44142 14744 44214
rect 14818 44204 14828 44214
rect 14818 44202 26089 44204
rect 14818 44146 26014 44202
rect 14818 44142 14828 44146
rect 25992 44144 26014 44146
rect 26078 44146 26089 44202
rect 26078 44144 26088 44146
rect 17668 44006 17678 44078
rect 17752 44066 17762 44078
rect 25444 44066 25454 44068
rect 17752 44014 25454 44066
rect 25510 44066 25520 44068
rect 25510 44014 25544 44066
rect 17752 44010 25544 44014
rect 17752 44006 17762 44010
rect 20614 43864 20624 43936
rect 20698 43926 20708 43936
rect 20698 43870 24898 43926
rect 20698 43864 20708 43870
rect 24888 43856 24898 43870
rect 24974 43870 25008 43926
rect 24974 43856 24984 43870
rect 23576 43768 23628 43778
rect 23560 43696 23570 43768
rect 23644 43760 23654 43768
rect 23644 43754 24432 43760
rect 23644 43708 24350 43754
rect 23644 43696 23654 43708
rect 24340 43684 24350 43708
rect 24426 43684 24436 43754
rect 26518 43568 26574 43570
rect 26516 43562 26578 43568
rect 26508 43550 26518 43562
rect 23785 43546 26518 43550
rect 23780 43482 23790 43546
rect 23854 43490 26518 43546
rect 26592 43490 26602 43562
rect 23854 43488 26578 43490
rect 23854 43482 23864 43488
rect 200 17360 17400 17380
rect 200 17200 220 17360
rect 560 17200 17400 17360
rect 200 17180 17400 17200
rect 220 16980 4140 17000
rect 220 16820 240 16980
rect 580 16820 4140 16980
rect 220 16800 4140 16820
rect 17200 16380 17400 17180
rect 13334 15026 14360 15040
rect 13334 14866 13354 15026
rect 13514 14866 14360 15026
rect 13334 14840 14360 14866
rect 7310 14400 7320 14580
rect 7480 14400 7490 14580
rect 9660 12280 9680 12460
rect 9860 12280 14360 12460
rect 9660 12260 14360 12280
rect 12540 12140 14240 12160
rect 12540 11980 12560 12140
rect 12740 11980 14240 12140
rect 12540 11960 14240 11980
rect 10180 11800 14360 11820
rect 810 11500 820 11720
rect 1160 11700 1170 11720
rect 1160 11500 3640 11700
rect 10180 11640 10200 11800
rect 10360 11640 14360 11800
rect 10180 11620 14360 11640
rect 12520 11240 14360 11260
rect 12520 11080 12540 11240
rect 12720 11080 14360 11240
rect 12520 11060 14360 11080
rect 810 10860 820 10880
rect 800 10700 820 10860
rect 810 10660 820 10700
rect 1160 10860 1170 10880
rect 1160 10700 14740 10860
rect 1160 10660 1170 10700
rect 2440 10460 7520 10480
rect 2440 10300 2460 10460
rect 2620 10300 7320 10460
rect 2440 10280 7320 10300
rect 7480 10280 7520 10460
rect 220 10100 6320 10120
rect 220 9940 240 10100
rect 580 9940 6320 10100
rect 220 9920 6320 9940
rect 6120 9600 6320 9920
rect 9400 7300 12748 7320
rect 9400 7120 12560 7300
rect 12726 7120 12748 7300
rect 1810 6000 1820 6200
rect 2020 6180 2940 6200
rect 2020 6020 2440 6180
rect 2640 6020 2940 6180
rect 2020 6000 2940 6020
rect 2180 5680 2200 5880
rect 2380 5680 2940 5880
rect 820 2260 840 2460
rect 830 2240 840 2260
rect 1180 2260 3040 2460
rect 1180 2240 1190 2260
<< via1 >>
rect 5906 44626 5972 44690
rect 27660 44626 27724 44684
rect 8846 44466 8920 44538
rect 27126 44476 27190 44534
rect 11794 44308 11868 44380
rect 26558 44318 26622 44376
rect 14744 44142 14818 44214
rect 26014 44144 26078 44202
rect 17678 44006 17752 44078
rect 25454 44014 25510 44068
rect 20624 43864 20698 43936
rect 24898 43856 24974 43926
rect 23570 43696 23644 43768
rect 24350 43684 24426 43754
rect 23790 43482 23854 43546
rect 26518 43490 26592 43562
rect 220 17200 560 17360
rect 240 16820 580 16980
rect 13354 14866 13514 15026
rect 7320 14400 7480 14580
rect 9680 12280 9860 12460
rect 12560 11980 12740 12140
rect 820 11500 1160 11720
rect 10200 11640 10360 11800
rect 12540 11080 12720 11240
rect 820 10660 1160 10880
rect 2460 10300 2620 10460
rect 7320 10280 7480 10460
rect 240 9940 580 10100
rect 12560 7120 12726 7300
rect 1820 6000 2020 6200
rect 2440 6020 2640 6180
rect 2200 5680 2380 5880
rect 840 2240 1180 2460
<< metal2 >>
rect 24332 44894 24424 44904
rect 23792 44832 23884 44842
rect 23789 44756 23792 44797
rect 24332 44808 24424 44818
rect 24888 44854 24980 44864
rect 24340 44800 24410 44808
rect 23789 44746 23884 44756
rect 23789 44738 23860 44746
rect 5910 44700 5966 44720
rect 5906 44690 5972 44700
rect 5906 44616 5972 44626
rect 5910 43324 5966 44616
rect 8854 44548 8910 44570
rect 8846 44538 8920 44548
rect 8846 44456 8920 44466
rect 8854 43306 8910 44456
rect 11794 44380 11868 44390
rect 11794 44298 11868 44308
rect 11798 43276 11854 44298
rect 14742 44224 14798 44230
rect 14742 44214 14818 44224
rect 14742 44142 14744 44214
rect 14742 44132 14818 44142
rect 14742 43214 14798 44132
rect 17678 44078 17752 44088
rect 17678 43996 17752 44006
rect 17686 43312 17742 43996
rect 20624 43936 20698 43946
rect 20624 43854 20698 43864
rect 20630 43260 20686 43854
rect 23570 43768 23644 43778
rect 23570 43686 23644 43696
rect 23574 43274 23630 43686
rect 23789 43556 23851 44738
rect 24350 43764 24410 44800
rect 24888 44768 24980 44778
rect 25446 44844 25538 44854
rect 24896 44760 24962 44768
rect 24902 43936 24962 44760
rect 25446 44758 25538 44768
rect 25454 44068 25514 44758
rect 27654 44696 27728 44706
rect 27654 44602 27728 44612
rect 27120 44546 27194 44556
rect 27120 44452 27194 44462
rect 26552 44388 26626 44398
rect 26552 44294 26626 44304
rect 28367 44276 28509 44314
rect 26008 44214 26082 44224
rect 26008 44120 26082 44130
rect 28367 44182 28382 44276
rect 28492 44182 28509 44276
rect 25510 44014 25514 44068
rect 25454 44006 25514 44014
rect 25454 44004 25510 44006
rect 24898 43926 24974 43936
rect 24898 43846 24974 43856
rect 24350 43754 24426 43764
rect 24350 43674 24426 43684
rect 26518 43562 26592 43572
rect 23789 43546 23854 43556
rect 23789 43488 23790 43546
rect 23790 43472 23854 43482
rect 26518 43480 26592 43490
rect 26518 43300 26574 43480
rect 28367 31194 28509 44182
rect 28367 31100 28390 31194
rect 28500 31100 28509 31194
rect 28367 31063 28509 31100
rect 9680 19160 9860 19170
rect 9660 18980 9680 19160
rect 220 17360 560 17370
rect 220 17190 560 17200
rect 240 16980 580 16990
rect 240 16810 580 16820
rect 7300 14580 7500 14600
rect 7300 14400 7320 14580
rect 7480 14400 7500 14580
rect 820 11720 1160 11730
rect 820 11490 1160 11500
rect 820 10880 1160 10890
rect 820 10650 1160 10660
rect 2440 10460 2640 10480
rect 2440 10300 2460 10460
rect 2620 10300 2640 10460
rect 240 10100 580 10110
rect 240 9930 580 9940
rect 1820 6200 2020 6210
rect 2440 6180 2640 10300
rect 7300 10460 7500 14400
rect 9660 12460 9860 18980
rect 9660 12280 9680 12460
rect 9660 12260 9860 12280
rect 10184 18680 10384 18700
rect 10184 18520 10200 18680
rect 10340 18520 10384 18680
rect 10184 11800 10384 18520
rect 10184 11640 10200 11800
rect 10360 11640 10384 11800
rect 10184 11620 10384 11640
rect 12540 18200 12740 18220
rect 12540 18040 12560 18200
rect 12540 12140 12740 18040
rect 12540 11980 12560 12140
rect 12540 11240 12740 11980
rect 12720 11080 12740 11240
rect 12540 11060 12740 11080
rect 13334 15026 13534 15040
rect 13334 14866 13354 15026
rect 13514 14866 13534 15026
rect 7300 10280 7320 10460
rect 7480 10280 7500 10460
rect 7320 10270 7480 10280
rect 2440 6010 2640 6020
rect 12548 7300 12748 7320
rect 12548 7120 12560 7300
rect 12726 7120 12748 7300
rect 840 2460 1180 2470
rect 840 2230 1180 2240
rect 1820 1570 2020 6000
rect 2200 5880 2380 5890
rect 2180 5680 2200 5880
rect 2180 1920 2380 5680
rect 11640 3000 11820 3010
rect 2180 1720 2200 1920
rect 2200 1710 2380 1720
rect 11620 2800 11640 2980
rect 11620 1920 11820 2800
rect 11800 1720 11820 1920
rect 12548 2040 12748 7120
rect 12548 1860 12560 2040
rect 12726 1860 12748 2040
rect 12548 1854 12748 1860
rect 12560 1850 12726 1854
rect 11620 1710 11800 1720
rect 1820 1560 2040 1570
rect 1820 1360 1840 1560
rect 1840 1350 2040 1360
rect 13334 1270 13534 14866
rect 13334 1110 13356 1270
rect 13516 1110 13534 1270
rect 13334 1076 13534 1110
<< via2 >>
rect 23792 44756 23884 44832
rect 24332 44818 24424 44894
rect 24888 44778 24980 44854
rect 25446 44768 25538 44844
rect 27654 44684 27728 44696
rect 27654 44626 27660 44684
rect 27660 44626 27724 44684
rect 27724 44626 27728 44684
rect 27654 44612 27728 44626
rect 27120 44534 27194 44546
rect 27120 44476 27126 44534
rect 27126 44476 27190 44534
rect 27190 44476 27194 44534
rect 27120 44462 27194 44476
rect 26552 44376 26626 44388
rect 26552 44318 26558 44376
rect 26558 44318 26622 44376
rect 26622 44318 26626 44376
rect 26552 44304 26626 44318
rect 26008 44202 26082 44214
rect 26008 44144 26014 44202
rect 26014 44144 26078 44202
rect 26078 44144 26082 44202
rect 26008 44130 26082 44144
rect 28382 44182 28492 44276
rect 28390 31100 28500 31194
rect 9680 18980 9860 19160
rect 220 17200 560 17360
rect 240 16820 580 16980
rect 820 11500 1160 11720
rect 820 10660 1160 10880
rect 240 9940 580 10100
rect 10200 18520 10340 18680
rect 12560 18040 12740 18200
rect 840 2240 1180 2460
rect 2200 1720 2380 1920
rect 11640 2800 11820 3000
rect 11620 1720 11800 1920
rect 12560 1860 12726 2040
rect 1840 1360 2040 1560
rect 13356 1110 13516 1270
<< metal3 >>
rect 24322 44894 24434 44899
rect 23782 44832 23894 44837
rect 23782 44756 23792 44832
rect 23884 44756 23894 44832
rect 24322 44818 24332 44894
rect 24424 44818 24434 44894
rect 24322 44813 24434 44818
rect 24878 44854 24990 44859
rect 24878 44778 24888 44854
rect 24980 44778 24990 44854
rect 24878 44773 24990 44778
rect 25436 44844 25548 44849
rect 25436 44768 25446 44844
rect 25538 44768 25548 44844
rect 25436 44763 25548 44768
rect 23782 44751 23894 44756
rect 27642 44696 27746 44714
rect 27642 44612 27654 44696
rect 27728 44612 27746 44696
rect 27642 44602 27746 44612
rect 27108 44546 27212 44564
rect 27108 44462 27120 44546
rect 27194 44462 27212 44546
rect 27108 44452 27212 44462
rect 26540 44388 26644 44406
rect 2910 44360 2920 44380
rect 2900 44200 2920 44360
rect 3100 44360 3110 44380
rect 3100 44340 15120 44360
rect 3100 44200 14920 44340
rect 2900 44160 14920 44200
rect 15100 44160 15120 44340
rect 26540 44304 26552 44388
rect 26626 44304 26644 44388
rect 26540 44294 26644 44304
rect 28180 44308 28509 44314
rect 25996 44214 26100 44232
rect 25996 44130 26008 44214
rect 26082 44130 26100 44214
rect 28180 44164 28194 44308
rect 28184 44162 28194 44164
rect 28304 44276 28509 44308
rect 28304 44182 28382 44276
rect 28492 44182 28509 44276
rect 28304 44172 28509 44182
rect 28304 44164 28322 44172
rect 28304 44162 28314 44164
rect 25996 44120 26100 44130
rect 3640 43980 28860 44000
rect 3640 43820 3660 43980
rect 3800 43820 28720 43980
rect 3640 43800 28720 43820
rect 28840 43800 28860 43980
rect 18778 43512 28208 43528
rect 18778 43508 28092 43512
rect 18778 43414 18802 43508
rect 18912 43418 28092 43508
rect 28202 43418 28212 43512
rect 18912 43414 28208 43418
rect 18778 43408 28208 43414
rect 220 43260 8180 43280
rect 220 43060 260 43260
rect 580 43060 7960 43260
rect 8140 43060 8180 43260
rect 220 43040 8180 43060
rect 28086 38986 28096 39080
rect 28206 38986 28216 39080
rect 28054 31199 28496 31204
rect 28054 31194 28510 31199
rect 28054 31100 28390 31194
rect 28500 31100 28510 31194
rect 28054 31095 28510 31100
rect 28054 31084 28496 31095
rect 28072 23296 28852 23316
rect 28072 23204 28728 23296
rect 28832 23204 28852 23296
rect 28072 23196 28852 23204
rect 806 19332 816 19526
rect 1154 19516 1164 19526
rect 1154 19500 8900 19516
rect 1154 19360 8680 19500
rect 8820 19360 8900 19500
rect 1154 19332 8900 19360
rect 830 19324 8900 19332
rect 9670 19160 9870 19165
rect 2900 19140 9680 19160
rect 2890 18960 2900 19140
rect 3080 18980 9680 19140
rect 9860 18980 9870 19160
rect 3080 18975 9870 18980
rect 3080 18960 9860 18975
rect 3640 18680 10384 18700
rect 3640 18520 3660 18680
rect 3800 18520 10200 18680
rect 10340 18520 10384 18680
rect 3640 18500 10384 18520
rect 200 18205 12740 18220
rect 200 18200 12750 18205
rect 200 18040 240 18200
rect 580 18040 12560 18200
rect 12740 18040 12750 18200
rect 200 18035 12750 18040
rect 200 18020 12740 18035
rect 210 17360 570 17365
rect 210 17200 220 17360
rect 560 17200 570 17360
rect 210 17195 570 17200
rect 230 16980 590 16985
rect 230 16820 240 16980
rect 580 16820 590 16980
rect 230 16815 590 16820
rect 810 11720 1170 11725
rect 810 11500 820 11720
rect 1160 11500 1170 11720
rect 810 11495 1170 11500
rect 810 10880 1170 10885
rect 810 10660 820 10880
rect 1160 10660 1170 10880
rect 810 10655 1170 10660
rect 230 10100 590 10105
rect 230 9940 240 10100
rect 580 9940 590 10100
rect 230 9935 590 9940
rect 11630 3000 11830 3005
rect 11630 2980 11640 3000
rect 11620 2800 11640 2980
rect 11820 2980 11830 3000
rect 11820 2800 22640 2980
rect 11620 2780 22640 2800
rect 22820 2780 22840 2980
rect 830 2460 1190 2465
rect 830 2240 840 2460
rect 1180 2240 1190 2460
rect 830 2235 1190 2240
rect 12548 2040 26698 2054
rect 2190 1920 2390 1925
rect 11610 1920 11810 1925
rect 2180 1720 2200 1920
rect 2380 1720 11620 1920
rect 11800 1720 11820 1920
rect 12548 1860 12560 2040
rect 12726 1860 26500 2040
rect 26666 1860 26698 2040
rect 12548 1854 26698 1860
rect 2190 1715 2390 1720
rect 11610 1715 11810 1720
rect 1830 1560 2050 1565
rect 18750 1560 18760 1580
rect 1820 1360 1840 1560
rect 2040 1380 18760 1560
rect 18960 1380 18970 1580
rect 2040 1360 18960 1380
rect 1830 1355 2050 1360
rect 13334 1270 30526 1276
rect 13334 1110 13356 1270
rect 13516 1260 30526 1270
rect 13516 1110 30376 1260
rect 13334 1100 30376 1110
rect 30536 1100 30546 1260
rect 13334 1076 30526 1100
<< via3 >>
rect 23792 44756 23884 44832
rect 24332 44818 24424 44894
rect 24888 44778 24980 44854
rect 25446 44768 25538 44844
rect 27654 44612 27728 44696
rect 27120 44462 27194 44546
rect 2920 44200 3100 44380
rect 14920 44160 15100 44340
rect 26552 44304 26626 44388
rect 26008 44130 26082 44214
rect 28194 44162 28304 44308
rect 3660 43820 3800 43980
rect 28720 43800 28840 43980
rect 18802 43414 18912 43508
rect 28092 43418 28202 43512
rect 260 43060 580 43260
rect 7960 43060 8140 43260
rect 28096 38986 28206 39080
rect 28728 23204 28832 23296
rect 816 19332 1154 19526
rect 8680 19360 8820 19500
rect 2900 18960 3080 19140
rect 3660 18520 3800 18680
rect 240 18040 580 18200
rect 220 17200 560 17360
rect 240 16820 580 16980
rect 820 11500 1160 11720
rect 820 10660 1160 10880
rect 240 9940 580 10100
rect 22640 2780 22820 2980
rect 840 2240 1180 2460
rect 26500 1860 26666 2040
rect 18760 1380 18960 1580
rect 30376 1100 30536 1260
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 2919 44380 3101 44381
rect 2919 44360 2920 44380
rect 2900 44200 2920 44360
rect 3100 44200 3101 44380
rect 14966 44341 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 2900 44199 3101 44200
rect 14919 44340 15101 44341
rect 200 43260 600 44152
rect 200 43060 260 43260
rect 580 43060 600 43260
rect 200 18200 600 43060
rect 200 18040 240 18200
rect 580 18040 600 18200
rect 200 17360 600 18040
rect 200 17200 220 17360
rect 560 17200 600 17360
rect 200 16980 600 17200
rect 200 16820 240 16980
rect 580 16820 600 16980
rect 200 10100 600 16820
rect 200 9940 240 10100
rect 580 9940 600 10100
rect 200 1000 600 9940
rect 800 19526 1200 44152
rect 800 19332 816 19526
rect 1154 19332 1200 19526
rect 800 11720 1200 19332
rect 2900 19141 3100 44199
rect 14919 44160 14920 44340
rect 15100 44160 15101 44340
rect 14919 44159 15101 44160
rect 2899 19140 3100 19141
rect 2899 18960 2900 19140
rect 3080 18960 3100 19140
rect 3640 43980 3840 44000
rect 3640 43820 3660 43980
rect 3800 43820 3840 43980
rect 2899 18959 3081 18960
rect 3640 18680 3840 43820
rect 18830 43509 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44844 23858 45152
rect 24350 44906 24410 45152
rect 24340 44895 24410 44906
rect 24331 44894 24425 44895
rect 23798 44833 23860 44844
rect 23791 44832 23885 44833
rect 23791 44756 23792 44832
rect 23884 44756 23885 44832
rect 24331 44818 24332 44894
rect 24424 44818 24425 44894
rect 24902 44866 24962 45152
rect 24896 44855 24962 44866
rect 24331 44817 24425 44818
rect 24887 44854 24981 44855
rect 24887 44778 24888 44854
rect 24980 44778 24981 44854
rect 25454 44845 25514 45152
rect 24887 44777 24981 44778
rect 25445 44844 25539 44845
rect 25445 44768 25446 44844
rect 25538 44768 25539 44844
rect 25445 44767 25539 44768
rect 23791 44755 23885 44756
rect 23798 44740 23858 44755
rect 26006 44236 26066 45152
rect 26558 44410 26618 45152
rect 27110 44568 27170 45152
rect 27662 44714 27722 45152
rect 27642 44696 27746 44714
rect 27642 44612 27654 44696
rect 27728 44612 27746 44696
rect 27642 44602 27746 44612
rect 27110 44564 27188 44568
rect 27108 44546 27212 44564
rect 27108 44462 27120 44546
rect 27194 44462 27212 44546
rect 27108 44452 27212 44462
rect 26558 44406 26620 44410
rect 26540 44388 26644 44406
rect 26540 44304 26552 44388
rect 26626 44304 26644 44388
rect 28214 44309 28274 45152
rect 26540 44294 26644 44304
rect 28193 44308 28305 44309
rect 26006 44232 26076 44236
rect 25996 44214 26100 44232
rect 25996 44130 26008 44214
rect 26082 44130 26100 44214
rect 28193 44162 28194 44308
rect 28304 44162 28305 44308
rect 28193 44161 28305 44162
rect 25996 44120 26100 44130
rect 28766 43981 28826 45152
rect 29318 44952 29378 45152
rect 28719 43980 28841 43981
rect 28719 43800 28720 43980
rect 28840 43892 28841 43980
rect 28840 43800 28852 43892
rect 28719 43799 28852 43800
rect 28088 43512 28208 43528
rect 18801 43508 18913 43509
rect 18801 43414 18802 43508
rect 18912 43414 18913 43508
rect 18801 43413 18913 43414
rect 28088 43418 28092 43512
rect 28202 43418 28208 43512
rect 18830 43402 18890 43413
rect 7906 43260 8222 43278
rect 7906 43060 7960 43260
rect 8140 43060 8222 43260
rect 7906 42728 8222 43060
rect 28088 39080 28208 43418
rect 28088 38986 28096 39080
rect 28206 38986 28208 39080
rect 28088 38972 28208 38986
rect 28732 23297 28852 43799
rect 28727 23296 28852 23297
rect 28727 23204 28728 23296
rect 28832 23204 28852 23296
rect 28727 23203 28852 23204
rect 28732 23196 28852 23203
rect 8674 19500 8866 19876
rect 8674 19360 8680 19500
rect 8820 19360 8866 19500
rect 8674 19324 8866 19360
rect 3640 18520 3660 18680
rect 3800 18520 3840 18680
rect 3640 18500 3840 18520
rect 800 11500 820 11720
rect 1160 11500 1200 11720
rect 800 10880 1200 11500
rect 800 10660 820 10880
rect 1160 10660 1200 10880
rect 800 2460 1200 10660
rect 800 2240 840 2460
rect 1180 2240 1200 2460
rect 800 1000 1200 2240
rect 22634 2981 22814 2990
rect 22634 2980 22821 2981
rect 22634 2780 22640 2980
rect 22820 2780 22821 2980
rect 22634 2779 22821 2780
rect 18759 1580 18961 1581
rect 18759 1380 18760 1580
rect 18960 1380 18961 1580
rect 18759 1379 18961 1380
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 220
rect 14906 0 15086 260
rect 18770 0 18950 1379
rect 22634 0 22814 2779
rect 26498 2040 26678 2060
rect 26498 1860 26500 2040
rect 26666 1860 26678 2040
rect 26498 0 26678 1860
rect 30362 1260 30542 1276
rect 30362 1100 30376 1260
rect 30536 1100 30542 1260
rect 30362 0 30542 1100
<< comment >>
rect 4720 19800 4740 19820
use buffer  buffer_0 /foss/designs/tt09-temp-sensor-clock_divider/mag/temp-sensor/buffer/mag
timestamp 1707919911
transform 1 0 1840 0 1 3980
box 900 -1720 7760 5820
use clock_divider  clock_divider_0 /foss/designs/tt09-temp-sensor-clock_divider/mag/clock-divider/mag_gds
timestamp 1729294469
transform 1 0 4226 0 1 19324
box 514 496 24000 24000
use sensor  sensor_0 /foss/designs/tt09-temp-sensor-clock_divider/mag/temp-sensor/sensor/mag
timestamp 1699935153
transform 1 0 3920 0 1 14000
box -660 -2500 3580 3000
use sigma-delta  sigma-delta_0 /foss/designs/tt09-temp-sensor-clock_divider/mag/temp-sensor/sigma-delta_modulator/mag
timestamp 1729283034
transform 1 0 17340 0 1 11220
box -3180 -520 12140 5420
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 200 1000 600 44152 1 FreeSans 2 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
