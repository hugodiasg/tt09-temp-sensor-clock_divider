magic
tech sky130A
magscale 1 2
timestamp 1729272731
<< viali >>
rect 10057 23273 10091 23307
rect 17877 23273 17911 23307
rect 4813 23205 4847 23239
rect 7757 23205 7791 23239
rect 8125 23205 8159 23239
rect 10977 23205 11011 23239
rect 14933 23205 14967 23239
rect 15149 23205 15183 23239
rect 20453 23205 20487 23239
rect 1777 23137 1811 23171
rect 5825 23137 5859 23171
rect 7113 23137 7147 23171
rect 7297 23137 7331 23171
rect 10057 23137 10091 23171
rect 10517 23137 10551 23171
rect 13553 23137 13587 23171
rect 15577 23137 15611 23171
rect 15945 23137 15979 23171
rect 16957 23137 16991 23171
rect 17233 23137 17267 23171
rect 17417 23137 17451 23171
rect 17693 23137 17727 23171
rect 18705 23137 18739 23171
rect 18889 23137 18923 23171
rect 19441 23137 19475 23171
rect 19993 23137 20027 23171
rect 20177 23137 20211 23171
rect 20269 23137 20303 23171
rect 20637 23137 20671 23171
rect 20729 23137 20763 23171
rect 20913 23137 20947 23171
rect 22385 23137 22419 23171
rect 9689 23069 9723 23103
rect 10241 23069 10275 23103
rect 10333 23069 10367 23103
rect 11805 23069 11839 23103
rect 13829 23069 13863 23103
rect 15393 23069 15427 23103
rect 16313 23069 16347 23103
rect 19625 23069 19659 23103
rect 22569 23069 22603 23103
rect 15853 23001 15887 23035
rect 17509 23001 17543 23035
rect 1961 22933 1995 22967
rect 4905 22933 4939 22967
rect 6009 22933 6043 22967
rect 7113 22933 7147 22967
rect 10701 22933 10735 22967
rect 15117 22933 15151 22967
rect 15301 22933 15335 22967
rect 18705 22933 18739 22967
rect 20085 22933 20119 22967
rect 20821 22933 20855 22967
rect 4721 22729 4755 22763
rect 5089 22729 5123 22763
rect 5365 22729 5399 22763
rect 7573 22729 7607 22763
rect 7757 22729 7791 22763
rect 9045 22729 9079 22763
rect 9689 22729 9723 22763
rect 18337 22729 18371 22763
rect 18521 22729 18555 22763
rect 7297 22661 7331 22695
rect 9413 22661 9447 22695
rect 8125 22593 8159 22627
rect 8953 22593 8987 22627
rect 9137 22593 9171 22627
rect 9965 22593 9999 22627
rect 10241 22593 10275 22627
rect 11161 22593 11195 22627
rect 16129 22593 16163 22627
rect 19993 22593 20027 22627
rect 21005 22593 21039 22627
rect 21281 22593 21315 22627
rect 21465 22593 21499 22627
rect 21925 22593 21959 22627
rect 4997 22525 5031 22559
rect 5181 22525 5215 22559
rect 5917 22525 5951 22559
rect 6009 22525 6043 22559
rect 6377 22525 6411 22559
rect 6655 22525 6689 22559
rect 7021 22525 7055 22559
rect 7113 22525 7147 22559
rect 7849 22525 7883 22559
rect 7941 22525 7975 22559
rect 9045 22525 9079 22559
rect 9505 22525 9539 22559
rect 10517 22525 10551 22559
rect 11345 22525 11379 22559
rect 11529 22525 11563 22559
rect 12449 22525 12483 22559
rect 12725 22525 12759 22559
rect 14289 22525 14323 22559
rect 14749 22525 14783 22559
rect 15577 22525 15611 22559
rect 15669 22525 15703 22559
rect 15853 22525 15887 22559
rect 17417 22525 17451 22559
rect 17785 22525 17819 22559
rect 19073 22525 19107 22559
rect 19533 22525 19567 22559
rect 19901 22525 19935 22559
rect 20269 22525 20303 22559
rect 20453 22525 20487 22559
rect 20913 22525 20947 22559
rect 21557 22525 21591 22559
rect 22017 22525 22051 22559
rect 22201 22525 22235 22559
rect 18383 22491 18417 22525
rect 4537 22457 4571 22491
rect 4753 22457 4787 22491
rect 6285 22457 6319 22491
rect 6745 22457 6779 22491
rect 6929 22457 6963 22491
rect 7297 22457 7331 22491
rect 7389 22457 7423 22491
rect 8125 22457 8159 22491
rect 18153 22457 18187 22491
rect 18705 22457 18739 22491
rect 4905 22389 4939 22423
rect 6653 22389 6687 22423
rect 7599 22389 7633 22423
rect 12357 22389 12391 22423
rect 12541 22389 12575 22423
rect 12909 22389 12943 22423
rect 16037 22389 16071 22423
rect 22109 22389 22143 22423
rect 10149 22185 10183 22219
rect 11529 22185 11563 22219
rect 21925 22185 21959 22219
rect 22477 22185 22511 22219
rect 5917 22117 5951 22151
rect 6285 22117 6319 22151
rect 6745 22117 6779 22151
rect 11069 22117 11103 22151
rect 12725 22117 12759 22151
rect 13093 22117 13127 22151
rect 17601 22117 17635 22151
rect 17785 22117 17819 22151
rect 18521 22117 18555 22151
rect 19993 22117 20027 22151
rect 5273 22049 5307 22083
rect 6101 22049 6135 22083
rect 6653 22049 6687 22083
rect 6837 22049 6871 22083
rect 7021 22049 7055 22083
rect 7113 22049 7147 22083
rect 7205 22049 7239 22083
rect 7573 22049 7607 22083
rect 7757 22049 7791 22083
rect 8677 22049 8711 22083
rect 9321 22049 9355 22083
rect 9873 22049 9907 22083
rect 9965 22049 9999 22083
rect 10241 22049 10275 22083
rect 11713 22049 11747 22083
rect 12081 22049 12115 22083
rect 14473 22049 14507 22083
rect 14749 22049 14783 22083
rect 16129 22049 16163 22083
rect 16957 22049 16991 22083
rect 17509 22049 17543 22083
rect 17693 22049 17727 22083
rect 17969 22049 18003 22083
rect 18245 22049 18279 22083
rect 18337 22049 18371 22083
rect 18613 22049 18647 22083
rect 19073 22049 19107 22083
rect 19441 22049 19475 22083
rect 20177 22049 20211 22083
rect 20361 22049 20395 22083
rect 20453 22049 20487 22083
rect 21465 22049 21499 22083
rect 21557 22049 21591 22083
rect 21649 22049 21683 22083
rect 6377 21981 6411 22015
rect 7481 21981 7515 22015
rect 10149 21981 10183 22015
rect 10701 21981 10735 22015
rect 13645 21981 13679 22015
rect 16865 21981 16899 22015
rect 19901 21981 19935 22015
rect 21741 21981 21775 22015
rect 22385 21981 22419 22015
rect 22937 21981 22971 22015
rect 10517 21913 10551 21947
rect 11437 21913 11471 21947
rect 18521 21913 18555 21947
rect 22109 21913 22143 21947
rect 22569 21913 22603 21947
rect 5365 21845 5399 21879
rect 6469 21845 6503 21879
rect 7665 21845 7699 21879
rect 8217 21845 8251 21879
rect 17417 21845 17451 21879
rect 18153 21845 18187 21879
rect 20729 21845 20763 21879
rect 21281 21845 21315 21879
rect 6837 21641 6871 21675
rect 8217 21641 8251 21675
rect 17141 21641 17175 21675
rect 19533 21641 19567 21675
rect 19717 21641 19751 21675
rect 20913 21641 20947 21675
rect 21097 21641 21131 21675
rect 8125 21573 8159 21607
rect 10701 21573 10735 21607
rect 20085 21573 20119 21607
rect 21925 21573 21959 21607
rect 22385 21573 22419 21607
rect 7849 21505 7883 21539
rect 12449 21505 12483 21539
rect 14749 21505 14783 21539
rect 17693 21505 17727 21539
rect 17877 21505 17911 21539
rect 18705 21505 18739 21539
rect 19165 21505 19199 21539
rect 22109 21505 22143 21539
rect 7021 21437 7055 21471
rect 7297 21437 7331 21471
rect 7481 21437 7515 21471
rect 7941 21437 7975 21471
rect 8217 21437 8251 21471
rect 9597 21437 9631 21471
rect 10241 21437 10275 21471
rect 11161 21437 11195 21471
rect 12725 21437 12759 21471
rect 13829 21437 13863 21471
rect 14197 21437 14231 21471
rect 14565 21437 14599 21471
rect 15485 21437 15519 21471
rect 16221 21437 16255 21471
rect 16865 21437 16899 21471
rect 17141 21437 17175 21471
rect 17601 21437 17635 21471
rect 17785 21437 17819 21471
rect 18061 21437 18095 21471
rect 19073 21437 19107 21471
rect 19809 21437 19843 21471
rect 21189 21437 21223 21471
rect 21373 21437 21407 21471
rect 21465 21437 21499 21471
rect 7665 21369 7699 21403
rect 10425 21369 10459 21403
rect 12173 21369 12207 21403
rect 13553 21369 13587 21403
rect 14013 21369 14047 21403
rect 17049 21369 17083 21403
rect 19349 21369 19383 21403
rect 19565 21369 19599 21403
rect 19901 21369 19935 21403
rect 20085 21369 20119 21403
rect 20729 21369 20763 21403
rect 21557 21369 21591 21403
rect 7205 21301 7239 21335
rect 10885 21301 10919 21335
rect 13369 21301 13403 21335
rect 13645 21301 13679 21335
rect 14289 21301 14323 21335
rect 18245 21301 18279 21335
rect 20929 21301 20963 21335
rect 21287 21301 21321 21335
rect 22017 21301 22051 21335
rect 22569 21301 22603 21335
rect 6469 21097 6503 21131
rect 11069 21097 11103 21131
rect 12909 21097 12943 21131
rect 19257 21097 19291 21131
rect 9321 21029 9355 21063
rect 12449 21029 12483 21063
rect 13093 21029 13127 21063
rect 13309 21029 13343 21063
rect 4353 20961 4387 20995
rect 5457 20961 5491 20995
rect 5641 20961 5675 20995
rect 5825 20961 5859 20995
rect 6009 20961 6043 20995
rect 6101 20961 6135 20995
rect 6193 20961 6227 20995
rect 7297 20961 7331 20995
rect 7389 20961 7423 20995
rect 7573 20961 7607 20995
rect 7941 20961 7975 20995
rect 8493 20961 8527 20995
rect 10057 20961 10091 20995
rect 10333 20961 10367 20995
rect 10701 20961 10735 20995
rect 10977 20961 11011 20995
rect 11253 20961 11287 20995
rect 14197 20961 14231 20995
rect 14933 20961 14967 20995
rect 16405 20961 16439 20995
rect 17325 20961 17359 20995
rect 17509 20961 17543 20995
rect 19165 20961 19199 20995
rect 20821 20961 20855 20995
rect 21005 20961 21039 20995
rect 21281 20961 21315 20995
rect 21465 20961 21499 20995
rect 21741 20961 21775 20995
rect 4445 20893 4479 20927
rect 7665 20893 7699 20927
rect 8401 20893 8435 20927
rect 16313 20893 16347 20927
rect 17233 20893 17267 20927
rect 20913 20893 20947 20927
rect 4721 20825 4755 20859
rect 7573 20825 7607 20859
rect 8125 20825 8159 20859
rect 12725 20825 12759 20859
rect 13461 20825 13495 20859
rect 5641 20757 5675 20791
rect 7757 20757 7791 20791
rect 11437 20757 11471 20791
rect 13277 20757 13311 20791
rect 17509 20757 17543 20791
rect 20637 20757 20671 20791
rect 21925 20757 21959 20791
rect 6009 20553 6043 20587
rect 6377 20553 6411 20587
rect 12909 20553 12943 20587
rect 18705 20553 18739 20587
rect 5089 20485 5123 20519
rect 7297 20485 7331 20519
rect 4261 20417 4295 20451
rect 6101 20417 6135 20451
rect 7849 20417 7883 20451
rect 13185 20417 13219 20451
rect 18797 20417 18831 20451
rect 4169 20349 4203 20383
rect 4353 20349 4387 20383
rect 4445 20349 4479 20383
rect 4629 20349 4663 20383
rect 4997 20349 5031 20383
rect 5181 20349 5215 20383
rect 5273 20349 5307 20383
rect 5365 20349 5399 20383
rect 5549 20349 5583 20383
rect 6009 20349 6043 20383
rect 8033 20349 8067 20383
rect 8125 20349 8159 20383
rect 12725 20349 12759 20383
rect 12909 20349 12943 20383
rect 13093 20349 13127 20383
rect 13277 20349 13311 20383
rect 13737 20349 13771 20383
rect 13921 20349 13955 20383
rect 14381 20349 14415 20383
rect 14473 20349 14507 20383
rect 14657 20349 14691 20383
rect 14933 20349 14967 20383
rect 15761 20349 15795 20383
rect 16497 20349 16531 20383
rect 17601 20349 17635 20383
rect 17969 20349 18003 20383
rect 18705 20349 18739 20383
rect 20913 20349 20947 20383
rect 21097 20349 21131 20383
rect 21373 20349 21407 20383
rect 21649 20349 21683 20383
rect 21833 20349 21867 20383
rect 22117 20349 22151 20383
rect 22385 20349 22419 20383
rect 22569 20349 22603 20383
rect 4813 20281 4847 20315
rect 7021 20281 7055 20315
rect 13553 20281 13587 20315
rect 15209 20281 15243 20315
rect 21925 20281 21959 20315
rect 22477 20281 22511 20315
rect 5733 20213 5767 20247
rect 7481 20213 7515 20247
rect 7849 20213 7883 20247
rect 14197 20213 14231 20247
rect 17233 20213 17267 20247
rect 19073 20213 19107 20247
rect 21005 20213 21039 20247
rect 21189 20213 21223 20247
rect 22293 20213 22327 20247
rect 13093 20009 13127 20043
rect 5641 19941 5675 19975
rect 9413 19941 9447 19975
rect 11069 19941 11103 19975
rect 18705 19941 18739 19975
rect 19073 19941 19107 19975
rect 19257 19941 19291 19975
rect 4445 19873 4479 19907
rect 4629 19873 4663 19907
rect 5273 19873 5307 19907
rect 5549 19873 5583 19907
rect 5917 19873 5951 19907
rect 6837 19873 6871 19907
rect 8401 19873 8435 19907
rect 8769 19873 8803 19907
rect 10057 19873 10091 19907
rect 10977 19873 11011 19907
rect 11161 19873 11195 19907
rect 11437 19873 11471 19907
rect 12725 19873 12759 19907
rect 12817 19873 12851 19907
rect 13461 19873 13495 19907
rect 13737 19873 13771 19907
rect 13829 19873 13863 19907
rect 15761 19873 15795 19907
rect 15945 19873 15979 19907
rect 16405 19873 16439 19907
rect 16865 19873 16899 19907
rect 17509 19873 17543 19907
rect 17601 19873 17635 19907
rect 18245 19873 18279 19907
rect 18889 19873 18923 19907
rect 18981 19873 19015 19907
rect 19349 19873 19383 19907
rect 20913 19873 20947 19907
rect 21097 19873 21131 19907
rect 21925 19873 21959 19907
rect 4353 19805 4387 19839
rect 5135 19805 5169 19839
rect 9781 19805 9815 19839
rect 10701 19805 10735 19839
rect 12357 19805 12391 19839
rect 13553 19805 13587 19839
rect 14013 19805 14047 19839
rect 17233 19805 17267 19839
rect 17785 19805 17819 19839
rect 18061 19805 18095 19839
rect 4813 19737 4847 19771
rect 7113 19737 7147 19771
rect 15945 19737 15979 19771
rect 17693 19737 17727 19771
rect 4997 19669 5031 19703
rect 12541 19669 12575 19703
rect 18429 19669 18463 19703
rect 18705 19669 18739 19703
rect 19165 19669 19199 19703
rect 21097 19669 21131 19703
rect 21833 19669 21867 19703
rect 11437 19465 11471 19499
rect 19993 19465 20027 19499
rect 21373 19465 21407 19499
rect 22017 19465 22051 19499
rect 8217 19397 8251 19431
rect 15485 19397 15519 19431
rect 18153 19397 18187 19431
rect 19441 19397 19475 19431
rect 11253 19329 11287 19363
rect 11805 19329 11839 19363
rect 13921 19329 13955 19363
rect 14565 19329 14599 19363
rect 18981 19329 19015 19363
rect 20545 19329 20579 19363
rect 21465 19329 21499 19363
rect 4813 19261 4847 19295
rect 4997 19261 5031 19295
rect 5089 19261 5123 19295
rect 5365 19261 5399 19295
rect 5641 19261 5675 19295
rect 5825 19261 5859 19295
rect 6193 19261 6227 19295
rect 7113 19261 7147 19295
rect 7389 19261 7423 19295
rect 8769 19261 8803 19295
rect 8861 19261 8895 19295
rect 9045 19261 9079 19295
rect 10241 19261 10275 19295
rect 10425 19261 10459 19295
rect 11345 19261 11379 19295
rect 11621 19261 11655 19295
rect 12265 19261 12299 19295
rect 12357 19261 12391 19295
rect 12521 19261 12555 19295
rect 13829 19261 13863 19295
rect 15393 19261 15427 19295
rect 16313 19261 16347 19295
rect 17233 19261 17267 19295
rect 17601 19261 17635 19295
rect 19073 19261 19107 19295
rect 19901 19261 19935 19295
rect 20085 19261 20119 19295
rect 20269 19261 20303 19295
rect 20361 19261 20395 19295
rect 20637 19261 20671 19295
rect 20821 19261 20855 19295
rect 20913 19261 20947 19295
rect 21005 19261 21039 19295
rect 21361 19261 21395 19295
rect 22293 19261 22327 19295
rect 22569 19261 22603 19295
rect 6101 19193 6135 19227
rect 18521 19193 18555 19227
rect 19809 19193 19843 19227
rect 21281 19193 21315 19227
rect 22001 19193 22035 19227
rect 22201 19193 22235 19227
rect 22477 19193 22511 19227
rect 4813 19125 4847 19159
rect 5181 19125 5215 19159
rect 5549 19125 5583 19159
rect 8401 19125 8435 19159
rect 12725 19125 12759 19159
rect 16865 19125 16899 19159
rect 18061 19125 18095 19159
rect 18705 19125 18739 19159
rect 19349 19125 19383 19159
rect 20545 19125 20579 19159
rect 21741 19125 21775 19159
rect 21833 19125 21867 19159
rect 22391 19125 22425 19159
rect 8033 18921 8067 18955
rect 9321 18921 9355 18955
rect 19441 18921 19475 18955
rect 22477 18921 22511 18955
rect 8493 18853 8527 18887
rect 17601 18853 17635 18887
rect 17785 18853 17819 18887
rect 6193 18785 6227 18819
rect 6285 18785 6319 18819
rect 6653 18785 6687 18819
rect 6837 18785 6871 18819
rect 7849 18785 7883 18819
rect 8033 18785 8067 18819
rect 8217 18785 8251 18819
rect 8401 18785 8435 18819
rect 8585 18785 8619 18819
rect 9229 18785 9263 18819
rect 9505 18785 9539 18819
rect 9965 18785 9999 18819
rect 10425 18785 10459 18819
rect 10793 18785 10827 18819
rect 11437 18785 11471 18819
rect 12173 18785 12207 18819
rect 12357 18785 12391 18819
rect 13461 18785 13495 18819
rect 13645 18785 13679 18819
rect 14473 18785 14507 18819
rect 14841 18785 14875 18819
rect 15117 18785 15151 18819
rect 17509 18785 17543 18819
rect 18521 18785 18555 18819
rect 19073 18785 19107 18819
rect 19197 18785 19231 18819
rect 19533 18785 19567 18819
rect 19717 18785 19751 18819
rect 20821 18785 20855 18819
rect 21281 18785 21315 18819
rect 21373 18785 21407 18819
rect 22201 18785 22235 18819
rect 5825 18717 5859 18751
rect 5917 18717 5951 18751
rect 7665 18717 7699 18751
rect 11161 18717 11195 18751
rect 12081 18717 12115 18751
rect 15669 18717 15703 18751
rect 18613 18717 18647 18751
rect 18969 18717 19003 18751
rect 20729 18717 20763 18751
rect 21557 18717 21591 18751
rect 8769 18649 8803 18683
rect 17785 18649 17819 18683
rect 19533 18649 19567 18683
rect 6469 18581 6503 18615
rect 9505 18581 9539 18615
rect 12265 18581 12299 18615
rect 18797 18581 18831 18615
rect 20453 18581 20487 18615
rect 20637 18581 20671 18615
rect 21465 18581 21499 18615
rect 6377 18377 6411 18411
rect 11805 18377 11839 18411
rect 14841 18377 14875 18411
rect 21879 18377 21913 18411
rect 22017 18377 22051 18411
rect 21097 18309 21131 18343
rect 4169 18241 4203 18275
rect 4445 18241 4479 18275
rect 4997 18241 5031 18275
rect 6009 18241 6043 18275
rect 7021 18241 7055 18275
rect 7757 18241 7791 18275
rect 8033 18241 8067 18275
rect 8861 18241 8895 18275
rect 10885 18241 10919 18275
rect 11713 18241 11747 18275
rect 12541 18241 12575 18275
rect 15209 18241 15243 18275
rect 15485 18241 15519 18275
rect 16129 18241 16163 18275
rect 20545 18241 20579 18275
rect 20637 18241 20671 18275
rect 21005 18241 21039 18275
rect 22109 18241 22143 18275
rect 22385 18241 22419 18275
rect 4077 18173 4111 18207
rect 6101 18173 6135 18207
rect 6561 18173 6595 18207
rect 6745 18173 6779 18207
rect 7205 18173 7239 18207
rect 7665 18173 7699 18207
rect 8769 18173 8803 18207
rect 10333 18173 10367 18207
rect 10701 18173 10735 18207
rect 11989 18173 12023 18207
rect 12173 18173 12207 18207
rect 13553 18173 13587 18207
rect 13737 18173 13771 18207
rect 14013 18173 14047 18207
rect 14749 18173 14783 18207
rect 16037 18173 16071 18207
rect 16957 18173 16991 18207
rect 17325 18173 17359 18207
rect 20729 18173 20763 18207
rect 20821 18173 20855 18207
rect 21468 18173 21502 18207
rect 21741 18173 21775 18207
rect 22201 18173 22235 18207
rect 22293 18173 22327 18207
rect 22477 18173 22511 18207
rect 5825 18105 5859 18139
rect 6653 18105 6687 18139
rect 13369 18105 13403 18139
rect 7389 18037 7423 18071
rect 8401 18037 8435 18071
rect 10701 18037 10735 18071
rect 14197 18037 14231 18071
rect 16037 18037 16071 18071
rect 16313 18037 16347 18071
rect 20361 18037 20395 18071
rect 21465 18037 21499 18071
rect 21649 18037 21683 18071
rect 5181 17833 5215 17867
rect 8309 17833 8343 17867
rect 13369 17833 13403 17867
rect 13553 17833 13587 17867
rect 19631 17833 19665 17867
rect 20453 17833 20487 17867
rect 21373 17833 21407 17867
rect 21649 17833 21683 17867
rect 6929 17765 6963 17799
rect 8953 17765 8987 17799
rect 19533 17765 19567 17799
rect 22762 17765 22796 17799
rect 4813 17697 4847 17731
rect 5917 17697 5951 17731
rect 7941 17697 7975 17731
rect 8125 17697 8159 17731
rect 8217 17697 8251 17731
rect 8769 17697 8803 17731
rect 9137 17697 9171 17731
rect 9505 17697 9539 17731
rect 11161 17697 11195 17731
rect 11621 17697 11655 17731
rect 11805 17697 11839 17731
rect 13550 17697 13584 17731
rect 14289 17697 14323 17731
rect 16497 17697 16531 17731
rect 18705 17697 18739 17731
rect 18797 17697 18831 17731
rect 18981 17697 19015 17731
rect 19073 17697 19107 17731
rect 19165 17697 19199 17731
rect 19717 17697 19751 17731
rect 19809 17697 19843 17731
rect 20269 17697 20303 17731
rect 20821 17697 20855 17731
rect 21281 17697 21315 17731
rect 21465 17697 21499 17731
rect 4721 17629 4755 17663
rect 8677 17629 8711 17663
rect 10057 17629 10091 17663
rect 11069 17629 11103 17663
rect 14013 17629 14047 17663
rect 14197 17629 14231 17663
rect 16405 17629 16439 17663
rect 18613 17629 18647 17663
rect 20085 17629 20119 17663
rect 20637 17629 20671 17663
rect 20729 17629 20763 17663
rect 20913 17629 20947 17663
rect 23029 17629 23063 17663
rect 14657 17561 14691 17595
rect 7757 17493 7791 17527
rect 11529 17493 11563 17527
rect 11989 17493 12023 17527
rect 13921 17493 13955 17527
rect 16221 17493 16255 17527
rect 19441 17493 19475 17527
rect 21097 17493 21131 17527
rect 14565 17289 14599 17323
rect 16497 17289 16531 17323
rect 22661 17289 22695 17323
rect 17417 17221 17451 17255
rect 22569 17221 22603 17255
rect 8769 17153 8803 17187
rect 9689 17153 9723 17187
rect 11437 17153 11471 17187
rect 11805 17153 11839 17187
rect 12357 17153 12391 17187
rect 13921 17153 13955 17187
rect 14749 17153 14783 17187
rect 16037 17153 16071 17187
rect 17785 17153 17819 17187
rect 18981 17153 19015 17187
rect 23029 17153 23063 17187
rect 8861 17085 8895 17119
rect 10609 17085 10643 17119
rect 10793 17085 10827 17119
rect 11345 17085 11379 17119
rect 11989 17085 12023 17119
rect 14013 17085 14047 17119
rect 14473 17085 14507 17119
rect 15669 17085 15703 17119
rect 15853 17085 15887 17119
rect 16129 17085 16163 17119
rect 16681 17085 16715 17119
rect 16774 17085 16808 17119
rect 17187 17085 17221 17119
rect 17417 17085 17451 17119
rect 17601 17085 17635 17119
rect 17693 17085 17727 17119
rect 17877 17085 17911 17119
rect 18889 17085 18923 17119
rect 19717 17085 19751 17119
rect 19984 17085 20018 17119
rect 21189 17085 21223 17119
rect 21445 17085 21479 17119
rect 22845 17085 22879 17119
rect 10517 17017 10551 17051
rect 16957 17017 16991 17051
rect 17049 17017 17083 17051
rect 18153 17017 18187 17051
rect 18337 17017 18371 17051
rect 18521 17017 18555 17051
rect 9229 16949 9263 16983
rect 10793 16949 10827 16983
rect 11713 16949 11747 16983
rect 12265 16949 12299 16983
rect 14381 16949 14415 16983
rect 14749 16949 14783 16983
rect 15761 16949 15795 16983
rect 17325 16949 17359 16983
rect 19257 16949 19291 16983
rect 21097 16949 21131 16983
rect 10241 16745 10275 16779
rect 11529 16745 11563 16779
rect 12541 16745 12575 16779
rect 14749 16745 14783 16779
rect 22661 16745 22695 16779
rect 6101 16677 6135 16711
rect 9781 16677 9815 16711
rect 10977 16677 11011 16711
rect 21548 16677 21582 16711
rect 6009 16609 6043 16643
rect 6285 16609 6319 16643
rect 6561 16609 6595 16643
rect 6745 16609 6779 16643
rect 11529 16609 11563 16643
rect 12081 16609 12115 16643
rect 12600 16609 12634 16643
rect 13461 16609 13495 16643
rect 14013 16609 14047 16643
rect 14197 16609 14231 16643
rect 14473 16609 14507 16643
rect 15209 16609 15243 16643
rect 16681 16609 16715 16643
rect 17325 16609 17359 16643
rect 18889 16609 18923 16643
rect 11621 16541 11655 16575
rect 12909 16541 12943 16575
rect 13369 16541 13403 16575
rect 16773 16541 16807 16575
rect 17049 16541 17083 16575
rect 17509 16541 17543 16575
rect 18981 16541 19015 16575
rect 21281 16541 21315 16575
rect 10057 16473 10091 16507
rect 12725 16473 12759 16507
rect 6469 16405 6503 16439
rect 6653 16405 6687 16439
rect 12173 16405 12207 16439
rect 14657 16405 14691 16439
rect 15025 16405 15059 16439
rect 17141 16405 17175 16439
rect 19165 16405 19199 16439
rect 10057 16201 10091 16235
rect 21925 16201 21959 16235
rect 22937 16201 22971 16235
rect 5089 16133 5123 16167
rect 14473 16133 14507 16167
rect 16773 16133 16807 16167
rect 7297 16065 7331 16099
rect 7573 16065 7607 16099
rect 9597 16065 9631 16099
rect 11161 16065 11195 16099
rect 15025 16065 15059 16099
rect 16957 16065 16991 16099
rect 22477 16065 22511 16099
rect 4813 15997 4847 16031
rect 5089 15997 5123 16031
rect 5365 15997 5399 16031
rect 5457 15997 5491 16031
rect 5733 15997 5767 16031
rect 6009 15997 6043 16031
rect 6469 15997 6503 16031
rect 6745 15997 6779 16031
rect 7021 15997 7055 16031
rect 7665 15997 7699 16031
rect 9505 15997 9539 16031
rect 9965 15997 9999 16031
rect 11069 15997 11103 16031
rect 13921 15997 13955 16031
rect 14105 15997 14139 16031
rect 14381 15997 14415 16031
rect 14565 15997 14599 16031
rect 14657 15997 14691 16031
rect 14841 15997 14875 16031
rect 15117 15997 15151 16031
rect 15577 15997 15611 16031
rect 15853 15997 15887 16031
rect 16037 15997 16071 16031
rect 16497 15997 16531 16031
rect 16589 15997 16623 16031
rect 16773 15997 16807 16031
rect 17049 15997 17083 16031
rect 22293 15997 22327 16031
rect 22753 15997 22787 16031
rect 4905 15929 4939 15963
rect 5549 15929 5583 15963
rect 6101 15929 6135 15963
rect 6193 15929 6227 15963
rect 6311 15929 6345 15963
rect 6929 15929 6963 15963
rect 14013 15929 14047 15963
rect 22385 15929 22419 15963
rect 5181 15861 5215 15895
rect 5825 15861 5859 15895
rect 6561 15861 6595 15895
rect 9873 15861 9907 15895
rect 10425 15861 10459 15895
rect 11805 15861 11839 15895
rect 14197 15861 14231 15895
rect 15485 15861 15519 15895
rect 15669 15861 15703 15895
rect 17417 15861 17451 15895
rect 5825 15657 5859 15691
rect 6285 15657 6319 15691
rect 6837 15657 6871 15691
rect 19073 15657 19107 15691
rect 20085 15657 20119 15691
rect 4528 15589 4562 15623
rect 6653 15589 6687 15623
rect 17325 15589 17359 15623
rect 6009 15521 6043 15555
rect 6193 15521 6227 15555
rect 6469 15521 6503 15555
rect 6745 15521 6779 15555
rect 6929 15521 6963 15555
rect 7021 15521 7055 15555
rect 7205 15521 7239 15555
rect 7481 15521 7515 15555
rect 8033 15521 8067 15555
rect 8493 15521 8527 15555
rect 10149 15521 10183 15555
rect 11253 15521 11287 15555
rect 13185 15521 13219 15555
rect 13461 15521 13495 15555
rect 13553 15521 13587 15555
rect 13737 15521 13771 15555
rect 13829 15521 13863 15555
rect 14841 15521 14875 15555
rect 16405 15521 16439 15555
rect 16589 15521 16623 15555
rect 17509 15521 17543 15555
rect 19165 15521 19199 15555
rect 19993 15521 20027 15555
rect 21537 15521 21571 15555
rect 4261 15453 4295 15487
rect 7665 15453 7699 15487
rect 7849 15453 7883 15487
rect 8677 15453 8711 15487
rect 10057 15453 10091 15487
rect 10977 15453 11011 15487
rect 11069 15453 11103 15487
rect 14013 15453 14047 15487
rect 14749 15453 14783 15487
rect 16497 15453 16531 15487
rect 16865 15453 16899 15487
rect 16957 15453 16991 15487
rect 17049 15453 17083 15487
rect 17141 15453 17175 15487
rect 18981 15453 19015 15487
rect 20177 15453 20211 15487
rect 21281 15453 21315 15487
rect 13369 15385 13403 15419
rect 15209 15385 15243 15419
rect 17693 15385 17727 15419
rect 5641 15317 5675 15351
rect 7205 15317 7239 15351
rect 7297 15317 7331 15351
rect 8217 15317 8251 15351
rect 8309 15317 8343 15351
rect 9873 15317 9907 15351
rect 11437 15317 11471 15351
rect 16681 15317 16715 15351
rect 19533 15317 19567 15351
rect 19625 15317 19659 15351
rect 22661 15317 22695 15351
rect 6285 15113 6319 15147
rect 7389 15113 7423 15147
rect 8585 15113 8619 15147
rect 12081 15113 12115 15147
rect 13185 15113 13219 15147
rect 17785 15113 17819 15147
rect 20085 15113 20119 15147
rect 21373 15113 21407 15147
rect 6653 14977 6687 15011
rect 11621 14977 11655 15011
rect 12541 14977 12575 15011
rect 13001 14977 13035 15011
rect 14105 14977 14139 15011
rect 21465 14977 21499 15011
rect 21925 14977 21959 15011
rect 4905 14909 4939 14943
rect 5172 14909 5206 14943
rect 6837 14909 6871 14943
rect 6929 14909 6963 14943
rect 7205 14909 7239 14943
rect 7481 14909 7515 14943
rect 7757 14909 7791 14943
rect 8033 14909 8067 14943
rect 8217 14909 8251 14943
rect 8585 14909 8619 14943
rect 8953 14909 8987 14943
rect 9045 14909 9079 14943
rect 9229 14909 9263 14943
rect 11529 14909 11563 14943
rect 11989 14909 12023 14943
rect 12265 14909 12299 14943
rect 12357 14909 12391 14943
rect 12909 14909 12943 14943
rect 14197 14909 14231 14943
rect 16313 14909 16347 14943
rect 16580 14909 16614 14943
rect 17969 14909 18003 14943
rect 18061 14909 18095 14943
rect 18337 14909 18371 14943
rect 18705 14909 18739 14943
rect 20361 14909 20395 14943
rect 21189 14909 21223 14943
rect 21373 14909 21407 14943
rect 21833 14909 21867 14943
rect 22293 14909 22327 14943
rect 12817 14841 12851 14875
rect 13185 14841 13219 14875
rect 18950 14841 18984 14875
rect 22477 14841 22511 14875
rect 6929 14773 6963 14807
rect 7021 14773 7055 14807
rect 7573 14773 7607 14807
rect 8401 14773 8435 14807
rect 9137 14773 9171 14807
rect 11897 14773 11931 14807
rect 13553 14773 13587 14807
rect 17693 14773 17727 14807
rect 18521 14773 18555 14807
rect 20177 14773 20211 14807
rect 22109 14773 22143 14807
rect 5181 14569 5215 14603
rect 7113 14569 7147 14603
rect 9873 14569 9907 14603
rect 10793 14569 10827 14603
rect 12909 14569 12943 14603
rect 17693 14569 17727 14603
rect 18429 14569 18463 14603
rect 21097 14569 21131 14603
rect 22293 14569 22327 14603
rect 8401 14501 8435 14535
rect 10241 14501 10275 14535
rect 12173 14501 12207 14535
rect 12265 14501 12299 14535
rect 13001 14501 13035 14535
rect 19564 14501 19598 14535
rect 5089 14433 5123 14467
rect 6377 14433 6411 14467
rect 6561 14433 6595 14467
rect 6653 14433 6687 14467
rect 6745 14433 6779 14467
rect 6929 14433 6963 14467
rect 7205 14433 7239 14467
rect 7389 14439 7423 14473
rect 7484 14436 7518 14470
rect 7619 14433 7653 14467
rect 9876 14433 9910 14467
rect 10149 14433 10183 14467
rect 10517 14433 10551 14467
rect 11345 14433 11379 14467
rect 11989 14433 12023 14467
rect 12449 14433 12483 14467
rect 12550 14455 12584 14489
rect 13185 14433 13219 14467
rect 13921 14433 13955 14467
rect 14013 14433 14047 14467
rect 17601 14433 17635 14467
rect 19809 14433 19843 14467
rect 20821 14433 20855 14467
rect 21465 14433 21499 14467
rect 21925 14433 21959 14467
rect 22109 14433 22143 14467
rect 22385 14433 22419 14467
rect 22569 14433 22603 14467
rect 5365 14365 5399 14399
rect 6469 14365 6503 14399
rect 9413 14365 9447 14399
rect 10609 14365 10643 14399
rect 11437 14365 11471 14399
rect 11805 14365 11839 14399
rect 12633 14365 12667 14399
rect 13645 14365 13679 14399
rect 13737 14365 13771 14399
rect 17877 14365 17911 14399
rect 21100 14365 21134 14399
rect 21557 14365 21591 14399
rect 8125 14297 8159 14331
rect 9505 14297 9539 14331
rect 10977 14297 11011 14331
rect 12265 14297 12299 14331
rect 4721 14229 4755 14263
rect 7849 14229 7883 14263
rect 7941 14229 7975 14263
rect 10057 14229 10091 14263
rect 12725 14229 12759 14263
rect 12817 14229 12851 14263
rect 13461 14229 13495 14263
rect 13829 14229 13863 14263
rect 17233 14229 17267 14263
rect 20913 14229 20947 14263
rect 21833 14229 21867 14263
rect 22109 14229 22143 14263
rect 22477 14229 22511 14263
rect 5733 14025 5767 14059
rect 9597 14025 9631 14059
rect 11621 14025 11655 14059
rect 18153 14025 18187 14059
rect 19533 14025 19567 14059
rect 16681 13957 16715 13991
rect 19165 13957 19199 13991
rect 7665 13889 7699 13923
rect 8493 13889 8527 13923
rect 9505 13889 9539 13923
rect 11437 13889 11471 13923
rect 11805 13889 11839 13923
rect 13645 13889 13679 13923
rect 14289 13889 14323 13923
rect 15669 13889 15703 13923
rect 15853 13889 15887 13923
rect 20821 13889 20855 13923
rect 21189 13889 21223 13923
rect 21465 13889 21499 13923
rect 4353 13821 4387 13855
rect 7573 13821 7607 13855
rect 8401 13821 8435 13855
rect 8585 13821 8619 13855
rect 9413 13821 9447 13855
rect 11253 13821 11287 13855
rect 11529 13821 11563 13855
rect 13737 13821 13771 13855
rect 14381 13821 14415 13855
rect 16037 13821 16071 13855
rect 16497 13821 16531 13855
rect 16773 13821 16807 13855
rect 17029 13821 17063 13855
rect 18981 13821 19015 13855
rect 19441 13821 19475 13855
rect 20637 13821 20671 13855
rect 21097 13821 21131 13855
rect 4598 13753 4632 13787
rect 11069 13753 11103 13787
rect 20453 13753 20487 13787
rect 7941 13685 7975 13719
rect 9781 13685 9815 13719
rect 11805 13685 11839 13719
rect 14105 13685 14139 13719
rect 14749 13685 14783 13719
rect 15209 13685 15243 13719
rect 15577 13685 15611 13719
rect 16221 13685 16255 13719
rect 3893 13481 3927 13515
rect 4169 13481 4203 13515
rect 5641 13481 5675 13515
rect 6285 13481 6319 13515
rect 19533 13481 19567 13515
rect 20729 13481 20763 13515
rect 21439 13481 21473 13515
rect 4506 13413 4540 13447
rect 6193 13413 6227 13447
rect 16374 13413 16408 13447
rect 19901 13413 19935 13447
rect 21649 13413 21683 13447
rect 3709 13345 3743 13379
rect 3985 13345 4019 13379
rect 7941 13345 7975 13379
rect 8217 13345 8251 13379
rect 8401 13345 8435 13379
rect 8677 13345 8711 13379
rect 8769 13345 8803 13379
rect 10149 13345 10183 13379
rect 10241 13345 10275 13379
rect 10609 13345 10643 13379
rect 10793 13345 10827 13379
rect 11161 13345 11195 13379
rect 11253 13345 11287 13379
rect 11989 13345 12023 13379
rect 14565 13345 14599 13379
rect 14832 13345 14866 13379
rect 16129 13345 16163 13379
rect 19165 13345 19199 13379
rect 19349 13345 19383 13379
rect 19625 13345 19659 13379
rect 19993 13345 20027 13379
rect 20177 13345 20211 13379
rect 20545 13345 20579 13379
rect 20729 13345 20763 13379
rect 4261 13277 4295 13311
rect 6469 13277 6503 13311
rect 10057 13277 10091 13311
rect 10333 13277 10367 13311
rect 11069 13277 11103 13311
rect 11345 13277 11379 13311
rect 11897 13277 11931 13311
rect 19717 13277 19751 13311
rect 19901 13277 19935 13311
rect 5825 13209 5859 13243
rect 8079 13209 8113 13243
rect 8493 13209 8527 13243
rect 10701 13209 10735 13243
rect 12357 13209 12391 13243
rect 8309 13141 8343 13175
rect 9873 13141 9907 13175
rect 11529 13141 11563 13175
rect 15945 13141 15979 13175
rect 17509 13141 17543 13175
rect 19165 13141 19199 13175
rect 20085 13141 20119 13175
rect 21281 13141 21315 13175
rect 21465 13141 21499 13175
rect 10425 12937 10459 12971
rect 15209 12937 15243 12971
rect 16405 12937 16439 12971
rect 17601 12937 17635 12971
rect 14289 12869 14323 12903
rect 17785 12869 17819 12903
rect 21005 12869 21039 12903
rect 21741 12869 21775 12903
rect 13737 12801 13771 12835
rect 13829 12801 13863 12835
rect 15025 12801 15059 12835
rect 15853 12801 15887 12835
rect 17509 12801 17543 12835
rect 18797 12801 18831 12835
rect 19257 12801 19291 12835
rect 21373 12801 21407 12835
rect 22201 12801 22235 12835
rect 22661 12801 22695 12835
rect 4261 12733 4295 12767
rect 4537 12733 4571 12767
rect 6837 12733 6871 12767
rect 9514 12733 9548 12767
rect 9781 12733 9815 12767
rect 10609 12733 10643 12767
rect 10793 12733 10827 12767
rect 11713 12733 11747 12767
rect 14749 12733 14783 12767
rect 15393 12733 15427 12767
rect 15945 12733 15979 12767
rect 16037 12733 16071 12767
rect 17601 12733 17635 12767
rect 18889 12733 18923 12767
rect 20729 12733 20763 12767
rect 20821 12733 20855 12767
rect 21005 12733 21039 12767
rect 21465 12733 21499 12767
rect 22109 12733 22143 12767
rect 22753 12733 22787 12767
rect 4782 12665 4816 12699
rect 7104 12665 7138 12699
rect 14841 12665 14875 12699
rect 17325 12665 17359 12699
rect 4445 12597 4479 12631
rect 5917 12597 5951 12631
rect 8217 12597 8251 12631
rect 8401 12597 8435 12631
rect 11529 12597 11563 12631
rect 13921 12597 13955 12631
rect 14381 12597 14415 12631
rect 21097 12597 21131 12631
rect 22385 12597 22419 12631
rect 4813 12393 4847 12427
rect 5273 12393 5307 12427
rect 7481 12393 7515 12427
rect 8585 12393 8619 12427
rect 10793 12393 10827 12427
rect 12909 12393 12943 12427
rect 13645 12393 13679 12427
rect 21005 12393 21039 12427
rect 21833 12393 21867 12427
rect 5181 12325 5215 12359
rect 9680 12325 9714 12359
rect 12090 12325 12124 12359
rect 12817 12325 12851 12359
rect 13982 12325 14016 12359
rect 17325 12325 17359 12359
rect 21281 12325 21315 12359
rect 7665 12257 7699 12291
rect 7849 12257 7883 12291
rect 7941 12257 7975 12291
rect 8585 12257 8619 12291
rect 8769 12257 8803 12291
rect 13461 12257 13495 12291
rect 15393 12257 15427 12291
rect 16957 12257 16991 12291
rect 17233 12257 17267 12291
rect 17417 12257 17451 12291
rect 18153 12257 18187 12291
rect 18337 12257 18371 12291
rect 20821 12257 20855 12291
rect 21557 12257 21591 12291
rect 22017 12257 22051 12291
rect 22109 12257 22143 12291
rect 22293 12257 22327 12291
rect 22569 12257 22603 12291
rect 23029 12257 23063 12291
rect 5457 12189 5491 12223
rect 9413 12189 9447 12223
rect 12357 12189 12391 12223
rect 13093 12189 13127 12223
rect 13737 12189 13771 12223
rect 17095 12189 17129 12223
rect 21373 12189 21407 12223
rect 22753 12189 22787 12223
rect 21741 12121 21775 12155
rect 22845 12121 22879 12155
rect 10977 12053 11011 12087
rect 12449 12053 12483 12087
rect 15117 12053 15151 12087
rect 15209 12053 15243 12087
rect 18245 12053 18279 12087
rect 21281 12053 21315 12087
rect 22109 12053 22143 12087
rect 22385 12053 22419 12087
rect 5365 11849 5399 11883
rect 5733 11849 5767 11883
rect 6009 11849 6043 11883
rect 11529 11849 11563 11883
rect 13553 11849 13587 11883
rect 15117 11849 15151 11883
rect 19257 11849 19291 11883
rect 19993 11849 20027 11883
rect 20453 11849 20487 11883
rect 21005 11849 21039 11883
rect 15577 11781 15611 11815
rect 16221 11781 16255 11815
rect 19901 11781 19935 11815
rect 5181 11713 5215 11747
rect 6101 11713 6135 11747
rect 11161 11713 11195 11747
rect 15301 11713 15335 11747
rect 16405 11713 16439 11747
rect 18797 11713 18831 11747
rect 19441 11713 19475 11747
rect 20085 11713 20119 11747
rect 5457 11645 5491 11679
rect 5549 11645 5583 11679
rect 5641 11645 5675 11679
rect 6009 11645 6043 11679
rect 6285 11645 6319 11679
rect 7941 11645 7975 11679
rect 8125 11645 8159 11679
rect 11345 11645 11379 11679
rect 12173 11645 12207 11679
rect 14677 11645 14711 11679
rect 14933 11645 14967 11679
rect 15393 11645 15427 11679
rect 16037 11645 16071 11679
rect 16221 11645 16255 11679
rect 16575 11645 16609 11679
rect 17141 11647 17175 11681
rect 17233 11645 17267 11679
rect 18889 11645 18923 11679
rect 19533 11645 19567 11679
rect 20269 11645 20303 11679
rect 22385 11645 22419 11679
rect 15117 11577 15151 11611
rect 19993 11577 20027 11611
rect 22140 11577 22174 11611
rect 5181 11509 5215 11543
rect 5917 11509 5951 11543
rect 6469 11509 6503 11543
rect 8033 11509 8067 11543
rect 11989 11509 12023 11543
rect 16865 11509 16899 11543
rect 16957 11509 16991 11543
rect 6837 11305 6871 11339
rect 7313 11305 7347 11339
rect 9045 11305 9079 11339
rect 12909 11305 12943 11339
rect 20913 11305 20947 11339
rect 21097 11305 21131 11339
rect 22661 11305 22695 11339
rect 5825 11237 5859 11271
rect 6041 11237 6075 11271
rect 6561 11237 6595 11271
rect 7113 11237 7147 11271
rect 8585 11237 8619 11271
rect 11796 11237 11830 11271
rect 15117 11237 15151 11271
rect 5273 11169 5307 11203
rect 6285 11169 6319 11203
rect 6377 11169 6411 11203
rect 6653 11169 6687 11203
rect 6837 11169 6871 11203
rect 7665 11169 7699 11203
rect 7757 11169 7791 11203
rect 8033 11169 8067 11203
rect 8171 11169 8205 11203
rect 8493 11169 8527 11203
rect 8769 11169 8803 11203
rect 8861 11169 8895 11203
rect 10977 11169 11011 11203
rect 11253 11169 11287 11203
rect 11345 11169 11379 11203
rect 11437 11169 11471 11203
rect 14013 11169 14047 11203
rect 14197 11169 14231 11203
rect 14749 11169 14783 11203
rect 15209 11169 15243 11203
rect 16129 11169 16163 11203
rect 16313 11169 16347 11203
rect 16589 11169 16623 11203
rect 16773 11169 16807 11203
rect 18889 11169 18923 11203
rect 21537 11169 21571 11203
rect 5365 11101 5399 11135
rect 8309 11101 8343 11135
rect 11529 11101 11563 11135
rect 15025 11101 15059 11135
rect 18981 11101 19015 11135
rect 19257 11101 19291 11135
rect 21281 11101 21315 11135
rect 7941 11033 7975 11067
rect 11115 11033 11149 11067
rect 14887 11033 14921 11067
rect 20545 11033 20579 11067
rect 5549 10965 5583 10999
rect 6009 10965 6043 10999
rect 6193 10965 6227 10999
rect 6561 10965 6595 10999
rect 7297 10965 7331 10999
rect 7481 10965 7515 10999
rect 8401 10965 8435 10999
rect 8585 10965 8619 10999
rect 14197 10965 14231 10999
rect 16221 10965 16255 10999
rect 16773 10965 16807 10999
rect 20913 10965 20947 10999
rect 6285 10761 6319 10795
rect 8217 10761 8251 10795
rect 9045 10761 9079 10795
rect 11713 10761 11747 10795
rect 16405 10761 16439 10795
rect 17785 10761 17819 10795
rect 18245 10761 18279 10795
rect 20913 10761 20947 10795
rect 21097 10761 21131 10795
rect 21833 10761 21867 10795
rect 22293 10761 22327 10795
rect 7757 10693 7791 10727
rect 12173 10693 12207 10727
rect 17049 10693 17083 10727
rect 21649 10693 21683 10727
rect 5549 10625 5583 10659
rect 6561 10625 6595 10659
rect 8677 10625 8711 10659
rect 10425 10625 10459 10659
rect 10701 10625 10735 10659
rect 11621 10625 11655 10659
rect 11897 10625 11931 10659
rect 14105 10625 14139 10659
rect 16129 10625 16163 10659
rect 16773 10625 16807 10659
rect 17233 10625 17267 10659
rect 17877 10625 17911 10659
rect 6653 10557 6687 10591
rect 7481 10557 7515 10591
rect 7849 10557 7883 10591
rect 8033 10557 8067 10591
rect 8769 10557 8803 10591
rect 9229 10557 9263 10591
rect 9321 10557 9355 10591
rect 9597 10557 9631 10591
rect 9781 10557 9815 10591
rect 9873 10557 9907 10591
rect 10057 10557 10091 10591
rect 10333 10557 10367 10591
rect 10517 10557 10551 10591
rect 10793 10557 10827 10591
rect 11437 10557 11471 10591
rect 11989 10557 12023 10591
rect 12633 10557 12667 10591
rect 12817 10557 12851 10591
rect 14013 10557 14047 10591
rect 14289 10557 14323 10591
rect 14473 10557 14507 10591
rect 14657 10557 14691 10591
rect 14749 10557 14783 10591
rect 14933 10557 14967 10591
rect 16037 10557 16071 10591
rect 16681 10557 16715 10591
rect 17325 10557 17359 10591
rect 18061 10557 18095 10591
rect 20637 10557 20671 10591
rect 21281 10557 21315 10591
rect 21557 10557 21591 10591
rect 22109 10557 22143 10591
rect 5733 10489 5767 10523
rect 6193 10489 6227 10523
rect 7757 10489 7791 10523
rect 9045 10489 9079 10523
rect 9965 10489 9999 10523
rect 11713 10489 11747 10523
rect 17785 10489 17819 10523
rect 20913 10489 20947 10523
rect 21801 10489 21835 10523
rect 22017 10489 22051 10523
rect 5641 10421 5675 10455
rect 6101 10421 6135 10455
rect 6837 10421 6871 10455
rect 7573 10421 7607 10455
rect 8401 10421 8435 10455
rect 9505 10421 9539 10455
rect 9781 10421 9815 10455
rect 11161 10421 11195 10455
rect 11253 10421 11287 10455
rect 12817 10421 12851 10455
rect 13645 10421 13679 10455
rect 14841 10421 14875 10455
rect 17693 10421 17727 10455
rect 20729 10421 20763 10455
rect 21465 10421 21499 10455
rect 6469 10217 6503 10251
rect 8769 10217 8803 10251
rect 9413 10217 9447 10251
rect 14657 10217 14691 10251
rect 20821 10217 20855 10251
rect 5273 10149 5307 10183
rect 19380 10149 19414 10183
rect 19809 10149 19843 10183
rect 6285 10081 6319 10115
rect 8401 10081 8435 10115
rect 9045 10081 9079 10115
rect 10241 10081 10275 10115
rect 10977 10081 11011 10115
rect 11161 10081 11195 10115
rect 14197 10081 14231 10115
rect 14473 10081 14507 10115
rect 19625 10081 19659 10115
rect 19717 10081 19751 10115
rect 19901 10081 19935 10115
rect 21097 10081 21131 10115
rect 21557 10081 21591 10115
rect 21741 10081 21775 10115
rect 22109 10081 22143 10115
rect 5825 10013 5859 10047
rect 6193 10013 6227 10047
rect 8309 10013 8343 10047
rect 9137 10013 9171 10047
rect 10149 10013 10183 10047
rect 14289 10013 14323 10047
rect 20821 10013 20855 10047
rect 21833 10013 21867 10047
rect 5641 9945 5675 9979
rect 21925 9945 21959 9979
rect 5089 9877 5123 9911
rect 5273 9877 5307 9911
rect 10609 9877 10643 9911
rect 11161 9877 11195 9911
rect 14197 9877 14231 9911
rect 18245 9877 18279 9911
rect 21005 9877 21039 9911
rect 21373 9877 21407 9911
rect 22017 9877 22051 9911
rect 5733 9673 5767 9707
rect 6561 9673 6595 9707
rect 7297 9673 7331 9707
rect 12081 9673 12115 9707
rect 14105 9673 14139 9707
rect 14289 9673 14323 9707
rect 18337 9673 18371 9707
rect 19349 9673 19383 9707
rect 20177 9673 20211 9707
rect 21097 9673 21131 9707
rect 7113 9605 7147 9639
rect 11989 9605 12023 9639
rect 12541 9605 12575 9639
rect 18061 9605 18095 9639
rect 18521 9605 18555 9639
rect 20085 9605 20119 9639
rect 20453 9605 20487 9639
rect 20545 9605 20579 9639
rect 10885 9537 10919 9571
rect 11529 9537 11563 9571
rect 12173 9537 12207 9571
rect 13645 9537 13679 9571
rect 14657 9537 14691 9571
rect 20269 9537 20303 9571
rect 20361 9537 20395 9571
rect 22477 9537 22511 9571
rect 4077 9469 4111 9503
rect 4353 9469 4387 9503
rect 6009 9469 6043 9503
rect 6101 9469 6135 9503
rect 6745 9469 6779 9503
rect 7021 9469 7055 9503
rect 10977 9469 11011 9503
rect 11621 9469 11655 9503
rect 12357 9469 12391 9503
rect 13737 9469 13771 9503
rect 14565 9469 14599 9503
rect 16405 9469 16439 9503
rect 16589 9469 16623 9503
rect 17877 9469 17911 9503
rect 18797 9469 18831 9503
rect 19073 9469 19107 9503
rect 19441 9469 19475 9503
rect 19717 9469 19751 9503
rect 19993 9469 20027 9503
rect 20637 9469 20671 9503
rect 20729 9469 20763 9503
rect 22569 9469 22603 9503
rect 22753 9469 22787 9503
rect 4598 9401 4632 9435
rect 5825 9401 5859 9435
rect 6929 9401 6963 9435
rect 7481 9401 7515 9435
rect 12081 9401 12115 9435
rect 18153 9401 18187 9435
rect 18981 9401 19015 9435
rect 22232 9401 22266 9435
rect 22661 9401 22695 9435
rect 4261 9333 4295 9367
rect 6193 9333 6227 9367
rect 6377 9333 6411 9367
rect 7271 9333 7305 9367
rect 11345 9333 11379 9367
rect 16497 9333 16531 9367
rect 18353 9333 18387 9367
rect 19165 9333 19199 9367
rect 19533 9333 19567 9367
rect 19901 9333 19935 9367
rect 20913 9333 20947 9367
rect 5825 9129 5859 9163
rect 8049 9129 8083 9163
rect 14197 9129 14231 9163
rect 17509 9129 17543 9163
rect 17877 9129 17911 9163
rect 19625 9129 19659 9163
rect 20729 9129 20763 9163
rect 22661 9129 22695 9163
rect 7849 9061 7883 9095
rect 16396 9061 16430 9095
rect 18398 9061 18432 9095
rect 19809 9061 19843 9095
rect 20545 9061 20579 9095
rect 4261 8993 4295 9027
rect 4528 8993 4562 9027
rect 6938 8993 6972 9027
rect 7205 8993 7239 9027
rect 13185 8993 13219 9027
rect 13829 8993 13863 9027
rect 17785 8993 17819 9027
rect 18061 8993 18095 9027
rect 20177 8993 20211 9027
rect 20269 8993 20303 9027
rect 20361 8993 20395 9027
rect 20913 8993 20947 9027
rect 21537 8993 21571 9027
rect 22753 8993 22787 9027
rect 13921 8925 13955 8959
rect 16129 8925 16163 8959
rect 18153 8925 18187 8959
rect 20545 8925 20579 8959
rect 21281 8925 21315 8959
rect 22937 8857 22971 8891
rect 5641 8789 5675 8823
rect 8033 8789 8067 8823
rect 8217 8789 8251 8823
rect 13369 8789 13403 8823
rect 18061 8789 18095 8823
rect 19533 8789 19567 8823
rect 19809 8789 19843 8823
rect 4905 8585 4939 8619
rect 5365 8585 5399 8619
rect 6009 8585 6043 8619
rect 6285 8585 6319 8619
rect 15577 8585 15611 8619
rect 15853 8585 15887 8619
rect 17233 8585 17267 8619
rect 17693 8585 17727 8619
rect 20085 8585 20119 8619
rect 20637 8585 20671 8619
rect 21097 8585 21131 8619
rect 21373 8585 21407 8619
rect 22201 8585 22235 8619
rect 5457 8517 5491 8551
rect 7297 8517 7331 8551
rect 13553 8517 13587 8551
rect 14105 8517 14139 8551
rect 15669 8517 15703 8551
rect 16221 8517 16255 8551
rect 17049 8517 17083 8551
rect 17601 8517 17635 8551
rect 21281 8517 21315 8551
rect 5549 8449 5583 8483
rect 6193 8449 6227 8483
rect 7389 8449 7423 8483
rect 8217 8449 8251 8483
rect 10241 8449 10275 8483
rect 10425 8449 10459 8483
rect 11529 8449 11563 8483
rect 14657 8449 14691 8483
rect 16313 8449 16347 8483
rect 16865 8449 16899 8483
rect 17785 8449 17819 8483
rect 21557 8449 21591 8483
rect 21741 8449 21775 8483
rect 21833 8449 21867 8483
rect 4905 8381 4939 8415
rect 5181 8381 5215 8415
rect 5283 8359 5317 8393
rect 5917 8381 5951 8415
rect 6285 8381 6319 8415
rect 6469 8381 6503 8415
rect 7021 8381 7055 8415
rect 7573 8381 7607 8415
rect 7665 8381 7699 8415
rect 7757 8381 7791 8415
rect 8033 8381 8067 8415
rect 8585 8381 8619 8415
rect 8677 8381 8711 8415
rect 8953 8381 8987 8415
rect 10517 8381 10551 8415
rect 11069 8381 11103 8415
rect 11161 8381 11195 8415
rect 11713 8381 11747 8415
rect 11805 8381 11839 8415
rect 12541 8381 12575 8415
rect 13921 8381 13955 8415
rect 14473 8381 14507 8415
rect 14841 8381 14875 8415
rect 14933 8381 14967 8415
rect 15117 8381 15151 8415
rect 15209 8381 15243 8415
rect 15393 8381 15427 8415
rect 16497 8381 16531 8415
rect 16589 8381 16623 8415
rect 17509 8381 17543 8415
rect 18705 8381 18739 8415
rect 18961 8381 18995 8415
rect 20361 8381 20395 8415
rect 20453 8381 20487 8415
rect 20637 8381 20671 8415
rect 20729 8381 20763 8415
rect 21649 8381 21683 8415
rect 22477 8381 22511 8415
rect 6193 8313 6227 8347
rect 7297 8313 7331 8347
rect 7389 8313 7423 8347
rect 8401 8313 8435 8347
rect 8769 8313 8803 8347
rect 10793 8313 10827 8347
rect 13829 8313 13863 8347
rect 14657 8313 14691 8347
rect 17417 8313 17451 8347
rect 22169 8313 22203 8347
rect 22385 8313 22419 8347
rect 5089 8245 5123 8279
rect 7113 8245 7147 8279
rect 7849 8245 7883 8279
rect 10241 8245 10275 8279
rect 10977 8245 11011 8279
rect 11345 8245 11379 8279
rect 11529 8245 11563 8279
rect 12725 8245 12759 8279
rect 13737 8245 13771 8279
rect 14381 8245 14415 8279
rect 15853 8245 15887 8279
rect 16681 8245 16715 8279
rect 17207 8245 17241 8279
rect 21097 8245 21131 8279
rect 22017 8245 22051 8279
rect 22661 8245 22695 8279
rect 7757 8041 7791 8075
rect 7849 8041 7883 8075
rect 10041 8041 10075 8075
rect 10977 8041 11011 8075
rect 12541 8041 12575 8075
rect 14197 8041 14231 8075
rect 15761 8041 15795 8075
rect 17509 8041 17543 8075
rect 21465 8041 21499 8075
rect 6644 7973 6678 8007
rect 9505 7973 9539 8007
rect 10241 7973 10275 8007
rect 10701 7973 10735 8007
rect 13062 7973 13096 8007
rect 14473 7973 14507 8007
rect 15945 7973 15979 8007
rect 17877 7973 17911 8007
rect 6377 7905 6411 7939
rect 8962 7905 8996 7939
rect 9229 7905 9263 7939
rect 9321 7905 9355 7939
rect 10517 7905 10551 7939
rect 10790 7927 10824 7961
rect 12090 7905 12124 7939
rect 12449 7905 12483 7939
rect 12725 7905 12759 7939
rect 12817 7905 12851 7939
rect 14933 7905 14967 7939
rect 15025 7905 15059 7939
rect 15209 7905 15243 7939
rect 15669 7905 15703 7939
rect 16129 7905 16163 7939
rect 16396 7905 16430 7939
rect 17601 7905 17635 7939
rect 17693 7905 17727 7939
rect 22578 7905 22612 7939
rect 22845 7905 22879 7939
rect 12357 7837 12391 7871
rect 17877 7837 17911 7871
rect 9873 7769 9907 7803
rect 14289 7769 14323 7803
rect 14841 7769 14875 7803
rect 10057 7701 10091 7735
rect 10333 7701 10367 7735
rect 12725 7701 12759 7735
rect 14473 7701 14507 7735
rect 15393 7701 15427 7735
rect 15945 7701 15979 7735
rect 7849 7497 7883 7531
rect 8769 7497 8803 7531
rect 9781 7497 9815 7531
rect 11713 7497 11747 7531
rect 12725 7497 12759 7531
rect 13185 7497 13219 7531
rect 13369 7497 13403 7531
rect 14933 7497 14967 7531
rect 16957 7497 16991 7531
rect 20453 7497 20487 7531
rect 22109 7497 22143 7531
rect 5733 7429 5767 7463
rect 7665 7429 7699 7463
rect 8493 7429 8527 7463
rect 9321 7429 9355 7463
rect 9965 7429 9999 7463
rect 10057 7429 10091 7463
rect 20085 7429 20119 7463
rect 20269 7429 20303 7463
rect 8217 7361 8251 7395
rect 8677 7361 8711 7395
rect 9413 7361 9447 7395
rect 12633 7361 12667 7395
rect 21557 7361 21591 7395
rect 7389 7293 7423 7327
rect 8401 7293 8435 7327
rect 8769 7293 8803 7327
rect 8953 7293 8987 7327
rect 9045 7293 9079 7327
rect 9137 7293 9171 7327
rect 11437 7293 11471 7327
rect 11529 7293 11563 7327
rect 11713 7293 11747 7327
rect 12817 7293 12851 7327
rect 12909 7293 12943 7327
rect 13553 7293 13587 7327
rect 15577 7293 15611 7327
rect 15844 7293 15878 7327
rect 19165 7293 19199 7327
rect 19809 7293 19843 7327
rect 20177 7293 20211 7327
rect 22201 7293 22235 7327
rect 22477 7293 22511 7327
rect 6009 7225 6043 7259
rect 7849 7225 7883 7259
rect 8677 7225 8711 7259
rect 9321 7225 9355 7259
rect 11170 7225 11204 7259
rect 13001 7225 13035 7259
rect 13820 7225 13854 7259
rect 20637 7225 20671 7259
rect 21741 7225 21775 7259
rect 5549 7157 5583 7191
rect 7573 7157 7607 7191
rect 9781 7157 9815 7191
rect 13201 7157 13235 7191
rect 19073 7157 19107 7191
rect 19901 7157 19935 7191
rect 19993 7157 20027 7191
rect 20427 7157 20461 7191
rect 21649 7157 21683 7191
rect 10793 6953 10827 6987
rect 11161 6953 11195 6987
rect 13921 6953 13955 6987
rect 14105 6953 14139 6987
rect 16313 6953 16347 6987
rect 18587 6953 18621 6987
rect 20453 6953 20487 6987
rect 21741 6953 21775 6987
rect 22293 6953 22327 6987
rect 22569 6953 22603 6987
rect 5273 6885 5307 6919
rect 6561 6885 6595 6919
rect 7726 6885 7760 6919
rect 9680 6885 9714 6919
rect 12808 6885 12842 6919
rect 18797 6885 18831 6919
rect 20269 6885 20303 6919
rect 4813 6817 4847 6851
rect 6101 6817 6135 6851
rect 6469 6817 6503 6851
rect 6745 6817 6779 6851
rect 7481 6817 7515 6851
rect 10977 6817 11011 6851
rect 14013 6817 14047 6851
rect 14197 6817 14231 6851
rect 16129 6817 16163 6851
rect 18153 6817 18187 6851
rect 19073 6817 19107 6851
rect 19257 6817 19291 6851
rect 19625 6817 19659 6851
rect 19901 6817 19935 6851
rect 20545 6817 20579 6851
rect 20729 6817 20763 6851
rect 20821 6817 20855 6851
rect 21373 6817 21407 6851
rect 22017 6817 22051 6851
rect 22109 6817 22143 6851
rect 22477 6817 22511 6851
rect 22569 6817 22603 6851
rect 22753 6817 22787 6851
rect 5825 6749 5859 6783
rect 6009 6749 6043 6783
rect 6193 6749 6227 6783
rect 6285 6749 6319 6783
rect 9413 6749 9447 6783
rect 12541 6749 12575 6783
rect 19441 6749 19475 6783
rect 21465 6749 21499 6783
rect 21833 6749 21867 6783
rect 5089 6681 5123 6715
rect 5641 6681 5675 6715
rect 18429 6681 18463 6715
rect 21005 6681 21039 6715
rect 4997 6613 5031 6647
rect 5273 6613 5307 6647
rect 6929 6613 6963 6647
rect 8861 6613 8895 6647
rect 18337 6613 18371 6647
rect 18613 6613 18647 6647
rect 18889 6613 18923 6647
rect 19809 6613 19843 6647
rect 20269 6613 20303 6647
rect 20637 6613 20671 6647
rect 21557 6613 21591 6647
rect 21925 6613 21959 6647
rect 6377 6409 6411 6443
rect 7021 6409 7055 6443
rect 20085 6409 20119 6443
rect 20913 6409 20947 6443
rect 21557 6341 21591 6375
rect 22661 6341 22695 6375
rect 7665 6273 7699 6307
rect 17693 6273 17727 6307
rect 21097 6273 21131 6307
rect 21189 6273 21223 6307
rect 4353 6205 4387 6239
rect 4813 6205 4847 6239
rect 4905 6205 4939 6239
rect 4997 6205 5031 6239
rect 5253 6205 5287 6239
rect 6745 6205 6779 6239
rect 7205 6205 7239 6239
rect 7297 6205 7331 6239
rect 17601 6205 17635 6239
rect 17785 6205 17819 6239
rect 17877 6205 17911 6239
rect 18061 6205 18095 6239
rect 18153 6205 18187 6239
rect 18245 6205 18279 6239
rect 18705 6205 18739 6239
rect 18961 6205 18995 6239
rect 20453 6205 20487 6239
rect 20545 6205 20579 6239
rect 20637 6205 20671 6239
rect 20821 6205 20855 6239
rect 21281 6205 21315 6239
rect 21373 6205 21407 6239
rect 21925 6205 21959 6239
rect 22385 6205 22419 6239
rect 22569 6205 22603 6239
rect 22845 6205 22879 6239
rect 4629 6137 4663 6171
rect 6469 6137 6503 6171
rect 6837 6137 6871 6171
rect 21741 6137 21775 6171
rect 22109 6137 22143 6171
rect 4537 6069 4571 6103
rect 4905 6069 4939 6103
rect 6653 6069 6687 6103
rect 7389 6069 7423 6103
rect 18521 6069 18555 6103
rect 20177 6069 20211 6103
rect 21833 6069 21867 6103
rect 22201 6069 22235 6103
rect 4261 5865 4295 5899
rect 7455 5865 7489 5899
rect 19441 5865 19475 5899
rect 21097 5865 21131 5899
rect 22845 5865 22879 5899
rect 7665 5797 7699 5831
rect 18328 5797 18362 5831
rect 19984 5797 20018 5831
rect 5385 5729 5419 5763
rect 5641 5729 5675 5763
rect 6081 5729 6115 5763
rect 18061 5729 18095 5763
rect 19717 5729 19751 5763
rect 21465 5729 21499 5763
rect 21732 5729 21766 5763
rect 5825 5661 5859 5695
rect 7297 5593 7331 5627
rect 7205 5525 7239 5559
rect 7481 5525 7515 5559
rect 4997 5321 5031 5355
rect 6469 5321 6503 5355
rect 18889 5321 18923 5355
rect 21373 5321 21407 5355
rect 21649 5321 21683 5355
rect 19993 5185 20027 5219
rect 4813 5117 4847 5151
rect 5089 5117 5123 5151
rect 18797 5117 18831 5151
rect 18981 5117 19015 5151
rect 21465 5117 21499 5151
rect 21649 5117 21683 5151
rect 5334 5049 5368 5083
rect 20260 5049 20294 5083
rect 5825 4777 5859 4811
rect 20269 4777 20303 4811
rect 6009 4641 6043 4675
rect 20453 4641 20487 4675
rect 6285 4573 6319 4607
rect 6193 4505 6227 4539
rect 22753 4097 22787 4131
rect 23029 4029 23063 4063
<< metal1 >>
rect 15930 23468 15936 23520
rect 15988 23508 15994 23520
rect 18414 23508 18420 23520
rect 15988 23480 18420 23508
rect 15988 23468 15994 23480
rect 18414 23468 18420 23480
rect 18472 23468 18478 23520
rect 552 23418 23368 23440
rect 552 23366 19022 23418
rect 19074 23366 19086 23418
rect 19138 23366 19150 23418
rect 19202 23366 19214 23418
rect 19266 23366 19278 23418
rect 19330 23366 23368 23418
rect 552 23344 23368 23366
rect 1670 23264 1676 23316
rect 1728 23264 1734 23316
rect 10045 23307 10103 23313
rect 10045 23273 10057 23307
rect 10091 23304 10103 23307
rect 11514 23304 11520 23316
rect 10091 23276 11520 23304
rect 10091 23273 10103 23276
rect 10045 23267 10103 23273
rect 11514 23264 11520 23276
rect 11572 23264 11578 23316
rect 17865 23307 17923 23313
rect 17865 23304 17877 23307
rect 16960 23276 17877 23304
rect 1688 23168 1716 23264
rect 4614 23196 4620 23248
rect 4672 23236 4678 23248
rect 4801 23239 4859 23245
rect 4801 23236 4813 23239
rect 4672 23208 4813 23236
rect 4672 23196 4678 23208
rect 4801 23205 4813 23208
rect 4847 23205 4859 23239
rect 4801 23199 4859 23205
rect 7558 23196 7564 23248
rect 7616 23236 7622 23248
rect 7745 23239 7803 23245
rect 7745 23236 7757 23239
rect 7616 23208 7757 23236
rect 7616 23196 7622 23208
rect 7745 23205 7757 23208
rect 7791 23205 7803 23239
rect 7745 23199 7803 23205
rect 8113 23239 8171 23245
rect 8113 23205 8125 23239
rect 8159 23236 8171 23239
rect 8159 23208 10456 23236
rect 8159 23205 8171 23208
rect 8113 23199 8171 23205
rect 1765 23171 1823 23177
rect 1765 23168 1777 23171
rect 1688 23140 1777 23168
rect 1765 23137 1777 23140
rect 1811 23137 1823 23171
rect 1765 23131 1823 23137
rect 5810 23128 5816 23180
rect 5868 23128 5874 23180
rect 7101 23171 7159 23177
rect 7101 23137 7113 23171
rect 7147 23168 7159 23171
rect 7190 23168 7196 23180
rect 7147 23140 7196 23168
rect 7147 23137 7159 23140
rect 7101 23131 7159 23137
rect 7190 23128 7196 23140
rect 7248 23128 7254 23180
rect 7285 23171 7343 23177
rect 7285 23137 7297 23171
rect 7331 23168 7343 23171
rect 7650 23168 7656 23180
rect 7331 23140 7656 23168
rect 7331 23137 7343 23140
rect 7285 23131 7343 23137
rect 7650 23128 7656 23140
rect 7708 23128 7714 23180
rect 5902 23060 5908 23112
rect 5960 23100 5966 23112
rect 8128 23100 8156 23199
rect 10045 23171 10103 23177
rect 10045 23137 10057 23171
rect 10091 23168 10103 23171
rect 10091 23140 10180 23168
rect 10091 23137 10103 23140
rect 10045 23131 10103 23137
rect 5960 23072 8156 23100
rect 5960 23060 5966 23072
rect 9674 23060 9680 23112
rect 9732 23060 9738 23112
rect 10152 23044 10180 23140
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23069 10287 23103
rect 10229 23063 10287 23069
rect 6638 23032 6644 23044
rect 6012 23004 6644 23032
rect 1949 22967 2007 22973
rect 1949 22933 1961 22967
rect 1995 22964 2007 22967
rect 4338 22964 4344 22976
rect 1995 22936 4344 22964
rect 1995 22933 2007 22936
rect 1949 22927 2007 22933
rect 4338 22924 4344 22936
rect 4396 22924 4402 22976
rect 4890 22924 4896 22976
rect 4948 22924 4954 22976
rect 6012 22973 6040 23004
rect 6638 22992 6644 23004
rect 6696 23032 6702 23044
rect 6696 23004 7512 23032
rect 6696 22992 6702 23004
rect 7484 22976 7512 23004
rect 10134 22992 10140 23044
rect 10192 22992 10198 23044
rect 5997 22967 6055 22973
rect 5997 22933 6009 22967
rect 6043 22933 6055 22967
rect 5997 22927 6055 22933
rect 7098 22924 7104 22976
rect 7156 22924 7162 22976
rect 7466 22924 7472 22976
rect 7524 22924 7530 22976
rect 9490 22924 9496 22976
rect 9548 22964 9554 22976
rect 10244 22964 10272 23063
rect 10318 23060 10324 23112
rect 10376 23060 10382 23112
rect 10428 23100 10456 23208
rect 10686 23196 10692 23248
rect 10744 23236 10750 23248
rect 10965 23239 11023 23245
rect 10965 23236 10977 23239
rect 10744 23208 10977 23236
rect 10744 23196 10750 23208
rect 10965 23205 10977 23208
rect 11011 23205 11023 23239
rect 10965 23199 11023 23205
rect 14366 23196 14372 23248
rect 14424 23236 14430 23248
rect 15194 23245 15200 23248
rect 14921 23239 14979 23245
rect 14921 23236 14933 23239
rect 14424 23208 14933 23236
rect 14424 23196 14430 23208
rect 14921 23205 14933 23208
rect 14967 23205 14979 23239
rect 14921 23199 14979 23205
rect 15137 23239 15200 23245
rect 15137 23205 15149 23239
rect 15183 23205 15200 23239
rect 15137 23199 15200 23205
rect 10502 23128 10508 23180
rect 10560 23128 10566 23180
rect 13446 23128 13452 23180
rect 13504 23168 13510 23180
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 13504 23140 13553 23168
rect 13504 23128 13510 23140
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 14936 23168 14964 23199
rect 15194 23196 15200 23199
rect 15252 23236 15258 23248
rect 15252 23208 15976 23236
rect 15252 23196 15258 23208
rect 15948 23180 15976 23208
rect 15565 23171 15623 23177
rect 15565 23168 15577 23171
rect 14936 23140 15577 23168
rect 13541 23131 13599 23137
rect 15565 23137 15577 23140
rect 15611 23137 15623 23171
rect 15565 23131 15623 23137
rect 15930 23128 15936 23180
rect 15988 23128 15994 23180
rect 16960 23177 16988 23276
rect 17865 23273 17877 23276
rect 17911 23304 17923 23307
rect 20898 23304 20904 23316
rect 17911 23276 20904 23304
rect 17911 23273 17923 23276
rect 17865 23267 17923 23273
rect 20898 23264 20904 23276
rect 20956 23264 20962 23316
rect 17034 23196 17040 23248
rect 17092 23236 17098 23248
rect 20441 23239 20499 23245
rect 17092 23208 17724 23236
rect 17092 23196 17098 23208
rect 16945 23171 17003 23177
rect 16945 23137 16957 23171
rect 16991 23137 17003 23171
rect 17221 23171 17279 23177
rect 17221 23168 17233 23171
rect 16945 23131 17003 23137
rect 17052 23140 17233 23168
rect 10428 23072 10548 23100
rect 10520 23032 10548 23072
rect 11790 23060 11796 23112
rect 11848 23060 11854 23112
rect 13817 23103 13875 23109
rect 13817 23069 13829 23103
rect 13863 23100 13875 23103
rect 14550 23100 14556 23112
rect 13863 23072 14556 23100
rect 13863 23069 13875 23072
rect 13817 23063 13875 23069
rect 14550 23060 14556 23072
rect 14608 23060 14614 23112
rect 15381 23103 15439 23109
rect 15381 23100 15393 23103
rect 15120 23072 15393 23100
rect 14918 23032 14924 23044
rect 10520 23004 14924 23032
rect 14918 22992 14924 23004
rect 14976 22992 14982 23044
rect 9548 22936 10272 22964
rect 10689 22967 10747 22973
rect 9548 22924 9554 22936
rect 10689 22933 10701 22967
rect 10735 22964 10747 22967
rect 11238 22964 11244 22976
rect 10735 22936 11244 22964
rect 10735 22933 10747 22936
rect 10689 22927 10747 22933
rect 11238 22924 11244 22936
rect 11296 22924 11302 22976
rect 14642 22924 14648 22976
rect 14700 22964 14706 22976
rect 15120 22973 15148 23072
rect 15381 23069 15393 23072
rect 15427 23100 15439 23103
rect 16298 23100 16304 23112
rect 15427 23072 16304 23100
rect 15427 23069 15439 23072
rect 15381 23063 15439 23069
rect 16298 23060 16304 23072
rect 16356 23060 16362 23112
rect 17052 23044 17080 23140
rect 17221 23137 17233 23140
rect 17267 23137 17279 23171
rect 17221 23131 17279 23137
rect 17405 23171 17463 23177
rect 17405 23137 17417 23171
rect 17451 23137 17463 23171
rect 17405 23131 17463 23137
rect 15841 23035 15899 23041
rect 15841 23001 15853 23035
rect 15887 23032 15899 23035
rect 17034 23032 17040 23044
rect 15887 23004 17040 23032
rect 15887 23001 15899 23004
rect 15841 22995 15899 23001
rect 17034 22992 17040 23004
rect 17092 22992 17098 23044
rect 15105 22967 15163 22973
rect 15105 22964 15117 22967
rect 14700 22936 15117 22964
rect 14700 22924 14706 22936
rect 15105 22933 15117 22936
rect 15151 22933 15163 22967
rect 15105 22927 15163 22933
rect 15289 22967 15347 22973
rect 15289 22933 15301 22967
rect 15335 22964 15347 22967
rect 16114 22964 16120 22976
rect 15335 22936 16120 22964
rect 15335 22933 15347 22936
rect 15289 22927 15347 22933
rect 16114 22924 16120 22936
rect 16172 22964 16178 22976
rect 17420 22964 17448 23131
rect 17494 23128 17500 23180
rect 17552 23128 17558 23180
rect 17696 23177 17724 23208
rect 18156 23208 20392 23236
rect 17681 23171 17739 23177
rect 17681 23137 17693 23171
rect 17727 23137 17739 23171
rect 17681 23131 17739 23137
rect 17512 23100 17540 23128
rect 18156 23100 18184 23208
rect 18690 23128 18696 23180
rect 18748 23128 18754 23180
rect 18877 23171 18935 23177
rect 18877 23137 18889 23171
rect 18923 23168 18935 23171
rect 19334 23168 19340 23180
rect 18923 23140 19340 23168
rect 18923 23137 18935 23140
rect 18877 23131 18935 23137
rect 19334 23128 19340 23140
rect 19392 23128 19398 23180
rect 19426 23128 19432 23180
rect 19484 23128 19490 23180
rect 19981 23171 20039 23177
rect 19981 23137 19993 23171
rect 20027 23137 20039 23171
rect 19981 23131 20039 23137
rect 20165 23171 20223 23177
rect 20165 23137 20177 23171
rect 20211 23168 20223 23171
rect 20257 23171 20315 23177
rect 20257 23168 20269 23171
rect 20211 23140 20269 23168
rect 20211 23137 20223 23140
rect 20165 23131 20223 23137
rect 20257 23137 20269 23140
rect 20303 23137 20315 23171
rect 20364 23168 20392 23208
rect 20441 23205 20453 23239
rect 20487 23236 20499 23239
rect 20530 23236 20536 23248
rect 20487 23208 20536 23236
rect 20487 23205 20499 23208
rect 20441 23199 20499 23205
rect 20530 23196 20536 23208
rect 20588 23236 20594 23248
rect 20588 23208 20944 23236
rect 20588 23196 20594 23208
rect 20625 23171 20683 23177
rect 20625 23168 20637 23171
rect 20364 23140 20637 23168
rect 20257 23131 20315 23137
rect 20625 23137 20637 23140
rect 20671 23168 20683 23171
rect 20714 23168 20720 23180
rect 20671 23140 20720 23168
rect 20671 23137 20683 23140
rect 20625 23131 20683 23137
rect 17512 23072 18184 23100
rect 18414 23060 18420 23112
rect 18472 23100 18478 23112
rect 19613 23103 19671 23109
rect 19613 23100 19625 23103
rect 18472 23072 19625 23100
rect 18472 23060 18478 23072
rect 19613 23069 19625 23072
rect 19659 23100 19671 23103
rect 19886 23100 19892 23112
rect 19659 23072 19892 23100
rect 19659 23069 19671 23072
rect 19613 23063 19671 23069
rect 19886 23060 19892 23072
rect 19944 23060 19950 23112
rect 19996 23100 20024 23131
rect 20714 23128 20720 23140
rect 20772 23128 20778 23180
rect 20916 23177 20944 23208
rect 20901 23171 20959 23177
rect 20901 23137 20913 23171
rect 20947 23137 20959 23171
rect 20901 23131 20959 23137
rect 22278 23128 22284 23180
rect 22336 23168 22342 23180
rect 22373 23171 22431 23177
rect 22373 23168 22385 23171
rect 22336 23140 22385 23168
rect 22336 23128 22342 23140
rect 22373 23137 22385 23140
rect 22419 23137 22431 23171
rect 22373 23131 22431 23137
rect 19996 23072 20852 23100
rect 17497 23035 17555 23041
rect 17497 23001 17509 23035
rect 17543 23032 17555 23035
rect 17543 23004 17816 23032
rect 17543 23001 17555 23004
rect 17497 22995 17555 23001
rect 17788 22976 17816 23004
rect 16172 22936 17448 22964
rect 16172 22924 16178 22936
rect 17770 22924 17776 22976
rect 17828 22924 17834 22976
rect 18693 22967 18751 22973
rect 18693 22933 18705 22967
rect 18739 22964 18751 22967
rect 19058 22964 19064 22976
rect 18739 22936 19064 22964
rect 18739 22933 18751 22936
rect 18693 22927 18751 22933
rect 19058 22924 19064 22936
rect 19116 22924 19122 22976
rect 19610 22924 19616 22976
rect 19668 22964 19674 22976
rect 20824 22973 20852 23072
rect 20990 23060 20996 23112
rect 21048 23100 21054 23112
rect 22557 23103 22615 23109
rect 22557 23100 22569 23103
rect 21048 23072 22569 23100
rect 21048 23060 21054 23072
rect 22557 23069 22569 23072
rect 22603 23069 22615 23103
rect 22557 23063 22615 23069
rect 20073 22967 20131 22973
rect 20073 22964 20085 22967
rect 19668 22936 20085 22964
rect 19668 22924 19674 22936
rect 20073 22933 20085 22936
rect 20119 22933 20131 22967
rect 20073 22927 20131 22933
rect 20809 22967 20867 22973
rect 20809 22933 20821 22967
rect 20855 22964 20867 22967
rect 21542 22964 21548 22976
rect 20855 22936 21548 22964
rect 20855 22933 20867 22936
rect 20809 22927 20867 22933
rect 21542 22924 21548 22936
rect 21600 22924 21606 22976
rect 552 22874 23368 22896
rect 552 22822 3662 22874
rect 3714 22822 3726 22874
rect 3778 22822 3790 22874
rect 3842 22822 3854 22874
rect 3906 22822 3918 22874
rect 3970 22822 23368 22874
rect 552 22800 23368 22822
rect 4709 22763 4767 22769
rect 4709 22729 4721 22763
rect 4755 22760 4767 22763
rect 5077 22763 5135 22769
rect 5077 22760 5089 22763
rect 4755 22732 5089 22760
rect 4755 22729 4767 22732
rect 4709 22723 4767 22729
rect 5077 22729 5089 22732
rect 5123 22729 5135 22763
rect 5077 22723 5135 22729
rect 5353 22763 5411 22769
rect 5353 22729 5365 22763
rect 5399 22760 5411 22763
rect 5810 22760 5816 22772
rect 5399 22732 5816 22760
rect 5399 22729 5411 22732
rect 5353 22723 5411 22729
rect 5092 22692 5120 22723
rect 5810 22720 5816 22732
rect 5868 22720 5874 22772
rect 7374 22760 7380 22772
rect 6932 22732 7380 22760
rect 5258 22692 5264 22704
rect 5092 22664 5264 22692
rect 5258 22652 5264 22664
rect 5316 22692 5322 22704
rect 5316 22664 6132 22692
rect 5316 22652 5322 22664
rect 6104 22624 6132 22664
rect 5000 22596 5948 22624
rect 4614 22556 4620 22568
rect 4540 22528 4620 22556
rect 4540 22497 4568 22528
rect 4614 22516 4620 22528
rect 4672 22556 4678 22568
rect 4890 22556 4896 22568
rect 4672 22528 4896 22556
rect 4672 22516 4678 22528
rect 4890 22516 4896 22528
rect 4948 22516 4954 22568
rect 5000 22565 5028 22596
rect 5920 22568 5948 22596
rect 6012 22596 6132 22624
rect 4985 22559 5043 22565
rect 4985 22525 4997 22559
rect 5031 22525 5043 22559
rect 4985 22519 5043 22525
rect 5169 22559 5227 22565
rect 5169 22525 5181 22559
rect 5215 22525 5227 22559
rect 5169 22519 5227 22525
rect 4525 22491 4583 22497
rect 4525 22457 4537 22491
rect 4571 22457 4583 22491
rect 4525 22451 4583 22457
rect 4741 22491 4799 22497
rect 4741 22457 4753 22491
rect 4787 22488 4799 22491
rect 5000 22488 5028 22519
rect 4787 22460 5028 22488
rect 5184 22488 5212 22519
rect 5902 22516 5908 22568
rect 5960 22516 5966 22568
rect 6012 22565 6040 22596
rect 5997 22559 6055 22565
rect 5997 22525 6009 22559
rect 6043 22525 6055 22559
rect 6178 22556 6184 22568
rect 5997 22519 6055 22525
rect 6104 22528 6184 22556
rect 6104 22488 6132 22528
rect 6178 22516 6184 22528
rect 6236 22556 6242 22568
rect 6365 22559 6423 22565
rect 6365 22556 6377 22559
rect 6236 22528 6377 22556
rect 6236 22516 6242 22528
rect 6365 22525 6377 22528
rect 6411 22525 6423 22559
rect 6638 22556 6644 22568
rect 6601 22528 6644 22556
rect 6365 22519 6423 22525
rect 6638 22516 6644 22528
rect 6696 22516 6702 22568
rect 6932 22556 6960 22732
rect 7374 22720 7380 22732
rect 7432 22760 7438 22772
rect 7561 22763 7619 22769
rect 7561 22760 7573 22763
rect 7432 22732 7573 22760
rect 7432 22720 7438 22732
rect 7561 22729 7573 22732
rect 7607 22729 7619 22763
rect 7561 22723 7619 22729
rect 7650 22720 7656 22772
rect 7708 22760 7714 22772
rect 7745 22763 7803 22769
rect 7745 22760 7757 22763
rect 7708 22732 7757 22760
rect 7708 22720 7714 22732
rect 7745 22729 7757 22732
rect 7791 22729 7803 22763
rect 7745 22723 7803 22729
rect 7190 22652 7196 22704
rect 7248 22692 7254 22704
rect 7285 22695 7343 22701
rect 7285 22692 7297 22695
rect 7248 22664 7297 22692
rect 7248 22652 7254 22664
rect 7285 22661 7297 22664
rect 7331 22692 7343 22695
rect 7331 22664 7604 22692
rect 7331 22661 7343 22664
rect 7285 22655 7343 22661
rect 7009 22559 7067 22565
rect 7009 22556 7021 22559
rect 6748 22528 7021 22556
rect 6748 22497 6776 22528
rect 7009 22525 7021 22528
rect 7055 22525 7067 22559
rect 7009 22519 7067 22525
rect 7101 22559 7159 22565
rect 7101 22525 7113 22559
rect 7147 22556 7159 22559
rect 7147 22528 7420 22556
rect 7147 22525 7159 22528
rect 7101 22519 7159 22525
rect 5184 22460 6132 22488
rect 6273 22491 6331 22497
rect 4787 22457 4799 22460
rect 4741 22451 4799 22457
rect 6273 22457 6285 22491
rect 6319 22488 6331 22491
rect 6733 22491 6791 22497
rect 6733 22488 6745 22491
rect 6319 22460 6745 22488
rect 6319 22457 6331 22460
rect 6273 22451 6331 22457
rect 6733 22457 6745 22460
rect 6779 22457 6791 22491
rect 6733 22451 6791 22457
rect 6917 22491 6975 22497
rect 6917 22457 6929 22491
rect 6963 22457 6975 22491
rect 6917 22451 6975 22457
rect 4890 22380 4896 22432
rect 4948 22380 4954 22432
rect 6638 22380 6644 22432
rect 6696 22380 6702 22432
rect 6932 22420 6960 22451
rect 7190 22448 7196 22500
rect 7248 22448 7254 22500
rect 7392 22497 7420 22528
rect 7285 22491 7343 22497
rect 7285 22457 7297 22491
rect 7331 22457 7343 22491
rect 7285 22451 7343 22457
rect 7377 22491 7435 22497
rect 7377 22457 7389 22491
rect 7423 22488 7435 22491
rect 7466 22488 7472 22500
rect 7423 22460 7472 22488
rect 7423 22457 7435 22460
rect 7377 22451 7435 22457
rect 7208 22420 7236 22448
rect 6932 22392 7236 22420
rect 7300 22420 7328 22451
rect 7466 22448 7472 22460
rect 7524 22448 7530 22500
rect 7576 22488 7604 22664
rect 7760 22556 7788 22723
rect 8478 22720 8484 22772
rect 8536 22760 8542 22772
rect 9033 22763 9091 22769
rect 9033 22760 9045 22763
rect 8536 22732 9045 22760
rect 8536 22720 8542 22732
rect 9033 22729 9045 22732
rect 9079 22729 9091 22763
rect 9033 22723 9091 22729
rect 9674 22720 9680 22772
rect 9732 22720 9738 22772
rect 10134 22720 10140 22772
rect 10192 22760 10198 22772
rect 10192 22732 10456 22760
rect 10192 22720 10198 22732
rect 9401 22695 9459 22701
rect 9401 22661 9413 22695
rect 9447 22692 9459 22695
rect 10318 22692 10324 22704
rect 9447 22664 10324 22692
rect 9447 22661 9459 22664
rect 9401 22655 9459 22661
rect 10318 22652 10324 22664
rect 10376 22652 10382 22704
rect 10428 22692 10456 22732
rect 16298 22720 16304 22772
rect 16356 22760 16362 22772
rect 18325 22763 18383 22769
rect 18325 22760 18337 22763
rect 16356 22732 18337 22760
rect 16356 22720 16362 22732
rect 18325 22729 18337 22732
rect 18371 22729 18383 22763
rect 18325 22723 18383 22729
rect 18509 22763 18567 22769
rect 18509 22729 18521 22763
rect 18555 22760 18567 22763
rect 18690 22760 18696 22772
rect 18555 22732 18696 22760
rect 18555 22729 18567 22732
rect 18509 22723 18567 22729
rect 18340 22692 18368 22723
rect 18690 22720 18696 22732
rect 18748 22720 18754 22772
rect 10428 22664 15884 22692
rect 18340 22664 20484 22692
rect 8110 22584 8116 22636
rect 8168 22584 8174 22636
rect 8941 22627 8999 22633
rect 8941 22593 8953 22627
rect 8987 22624 8999 22627
rect 9125 22627 9183 22633
rect 9125 22624 9137 22627
rect 8987 22596 9137 22624
rect 8987 22593 8999 22596
rect 8941 22587 8999 22593
rect 9125 22593 9137 22596
rect 9171 22624 9183 22627
rect 9953 22627 10011 22633
rect 9171 22596 9628 22624
rect 9171 22593 9183 22596
rect 9125 22587 9183 22593
rect 7837 22559 7895 22565
rect 7837 22556 7849 22559
rect 7760 22528 7849 22556
rect 7837 22525 7849 22528
rect 7883 22525 7895 22559
rect 7837 22519 7895 22525
rect 7926 22516 7932 22568
rect 7984 22516 7990 22568
rect 9030 22556 9036 22568
rect 8036 22528 9036 22556
rect 7944 22488 7972 22516
rect 8036 22500 8064 22528
rect 9030 22516 9036 22528
rect 9088 22516 9094 22568
rect 9490 22516 9496 22568
rect 9548 22516 9554 22568
rect 9600 22556 9628 22596
rect 9953 22593 9965 22627
rect 9999 22624 10011 22627
rect 10229 22627 10287 22633
rect 10229 22624 10241 22627
rect 9999 22596 10241 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 10229 22593 10241 22596
rect 10275 22593 10287 22627
rect 10229 22587 10287 22593
rect 10134 22556 10140 22568
rect 9600 22528 10140 22556
rect 10134 22516 10140 22528
rect 10192 22516 10198 22568
rect 10505 22559 10563 22565
rect 10505 22525 10517 22559
rect 10551 22556 10563 22559
rect 10888 22556 10916 22664
rect 11149 22627 11207 22633
rect 11149 22593 11161 22627
rect 11195 22624 11207 22627
rect 11422 22624 11428 22636
rect 11195 22596 11428 22624
rect 11195 22593 11207 22596
rect 11149 22587 11207 22593
rect 11422 22584 11428 22596
rect 11480 22624 11486 22636
rect 11480 22596 11560 22624
rect 11480 22584 11486 22596
rect 10551 22528 10916 22556
rect 10551 22525 10563 22528
rect 10505 22519 10563 22525
rect 11330 22516 11336 22568
rect 11388 22516 11394 22568
rect 11532 22565 11560 22596
rect 11974 22584 11980 22636
rect 12032 22624 12038 22636
rect 15856 22624 15884 22664
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 12032 22596 12756 22624
rect 12032 22584 12038 22596
rect 12728 22565 12756 22596
rect 15488 22596 15700 22624
rect 15856 22596 16129 22624
rect 11517 22559 11575 22565
rect 11517 22525 11529 22559
rect 11563 22525 11575 22559
rect 11517 22519 11575 22525
rect 12437 22559 12495 22565
rect 12437 22525 12449 22559
rect 12483 22525 12495 22559
rect 12437 22519 12495 22525
rect 12713 22559 12771 22565
rect 12713 22525 12725 22559
rect 12759 22525 12771 22559
rect 12713 22519 12771 22525
rect 14277 22559 14335 22565
rect 14277 22525 14289 22559
rect 14323 22556 14335 22559
rect 14366 22556 14372 22568
rect 14323 22528 14372 22556
rect 14323 22525 14335 22528
rect 14277 22519 14335 22525
rect 7576 22460 7972 22488
rect 8018 22448 8024 22500
rect 8076 22448 8082 22500
rect 8113 22491 8171 22497
rect 8113 22457 8125 22491
rect 8159 22488 8171 22491
rect 9508 22488 9536 22516
rect 8159 22460 9536 22488
rect 8159 22457 8171 22460
rect 8113 22451 8171 22457
rect 12452 22432 12480 22519
rect 14366 22516 14372 22528
rect 14424 22516 14430 22568
rect 14737 22559 14795 22565
rect 14737 22525 14749 22559
rect 14783 22525 14795 22559
rect 14737 22519 14795 22525
rect 13912 22500 13964 22506
rect 13912 22442 13964 22448
rect 7587 22423 7645 22429
rect 7587 22420 7599 22423
rect 7300 22392 7599 22420
rect 7587 22389 7599 22392
rect 7633 22420 7645 22423
rect 9490 22420 9496 22432
rect 7633 22392 9496 22420
rect 7633 22389 7645 22392
rect 7587 22383 7645 22389
rect 9490 22380 9496 22392
rect 9548 22380 9554 22432
rect 12345 22423 12403 22429
rect 12345 22389 12357 22423
rect 12391 22420 12403 22423
rect 12434 22420 12440 22432
rect 12391 22392 12440 22420
rect 12391 22389 12403 22392
rect 12345 22383 12403 22389
rect 12434 22380 12440 22392
rect 12492 22380 12498 22432
rect 12526 22380 12532 22432
rect 12584 22380 12590 22432
rect 12894 22380 12900 22432
rect 12952 22380 12958 22432
rect 14550 22380 14556 22432
rect 14608 22420 14614 22432
rect 14752 22420 14780 22519
rect 14918 22516 14924 22568
rect 14976 22556 14982 22568
rect 15378 22556 15384 22568
rect 14976 22528 15384 22556
rect 14976 22516 14982 22528
rect 15378 22516 15384 22528
rect 15436 22556 15442 22568
rect 15488 22556 15516 22596
rect 15436 22528 15516 22556
rect 15436 22516 15442 22528
rect 15562 22516 15568 22568
rect 15620 22516 15626 22568
rect 15672 22565 15700 22596
rect 16117 22593 16129 22596
rect 16163 22593 16175 22627
rect 18414 22624 18420 22636
rect 16117 22587 16175 22593
rect 18356 22596 18420 22624
rect 15657 22559 15715 22565
rect 15657 22525 15669 22559
rect 15703 22525 15715 22559
rect 15841 22559 15899 22565
rect 15841 22556 15853 22559
rect 15657 22519 15715 22525
rect 15764 22528 15853 22556
rect 15010 22448 15016 22500
rect 15068 22488 15074 22500
rect 15764 22488 15792 22528
rect 15841 22525 15853 22528
rect 15887 22556 15899 22559
rect 16132 22556 16160 22587
rect 17310 22556 17316 22568
rect 15887 22528 16068 22556
rect 16132 22528 17316 22556
rect 15887 22525 15899 22528
rect 15841 22519 15899 22525
rect 15068 22460 15792 22488
rect 16040 22488 16068 22528
rect 17310 22516 17316 22528
rect 17368 22516 17374 22568
rect 17402 22516 17408 22568
rect 17460 22516 17466 22568
rect 17770 22516 17776 22568
rect 17828 22516 17834 22568
rect 18356 22531 18384 22596
rect 18414 22584 18420 22596
rect 18472 22584 18478 22636
rect 19334 22584 19340 22636
rect 19392 22624 19398 22636
rect 19981 22627 20039 22633
rect 19981 22624 19993 22627
rect 19392 22596 19993 22624
rect 19392 22584 19398 22596
rect 19981 22593 19993 22596
rect 20027 22593 20039 22627
rect 19981 22587 20039 22593
rect 18356 22525 18429 22531
rect 16574 22488 16580 22500
rect 16040 22460 16580 22488
rect 15068 22448 15074 22460
rect 16574 22448 16580 22460
rect 16632 22448 16638 22500
rect 18141 22491 18199 22497
rect 18356 22494 18383 22525
rect 18141 22457 18153 22491
rect 18187 22457 18199 22491
rect 18371 22491 18383 22494
rect 18417 22491 18429 22525
rect 19058 22516 19064 22568
rect 19116 22516 19122 22568
rect 19518 22516 19524 22568
rect 19576 22516 19582 22568
rect 19886 22516 19892 22568
rect 19944 22516 19950 22568
rect 20456 22565 20484 22664
rect 20990 22584 20996 22636
rect 21048 22584 21054 22636
rect 21269 22627 21327 22633
rect 21269 22593 21281 22627
rect 21315 22624 21327 22627
rect 21450 22624 21456 22636
rect 21315 22596 21456 22624
rect 21315 22593 21327 22596
rect 21269 22587 21327 22593
rect 21450 22584 21456 22596
rect 21508 22584 21514 22636
rect 21910 22584 21916 22636
rect 21968 22584 21974 22636
rect 20257 22559 20315 22565
rect 20257 22525 20269 22559
rect 20303 22525 20315 22559
rect 20257 22519 20315 22525
rect 20441 22559 20499 22565
rect 20441 22525 20453 22559
rect 20487 22556 20499 22559
rect 20901 22559 20959 22565
rect 20901 22556 20913 22559
rect 20487 22528 20913 22556
rect 20487 22525 20499 22528
rect 20441 22519 20499 22525
rect 20901 22525 20913 22528
rect 20947 22525 20959 22559
rect 20901 22519 20959 22525
rect 18371 22485 18429 22491
rect 18141 22451 18199 22457
rect 15562 22420 15568 22432
rect 14608 22392 15568 22420
rect 14608 22380 14614 22392
rect 15562 22380 15568 22392
rect 15620 22380 15626 22432
rect 16025 22423 16083 22429
rect 16025 22389 16037 22423
rect 16071 22420 16083 22423
rect 17494 22420 17500 22432
rect 16071 22392 17500 22420
rect 16071 22389 16083 22392
rect 16025 22383 16083 22389
rect 17494 22380 17500 22392
rect 17552 22380 17558 22432
rect 17770 22380 17776 22432
rect 17828 22420 17834 22432
rect 18156 22420 18184 22451
rect 18598 22448 18604 22500
rect 18656 22488 18662 22500
rect 18693 22491 18751 22497
rect 18693 22488 18705 22491
rect 18656 22460 18705 22488
rect 18656 22448 18662 22460
rect 18693 22457 18705 22460
rect 18739 22457 18751 22491
rect 20272 22488 20300 22519
rect 21542 22516 21548 22568
rect 21600 22516 21606 22568
rect 22002 22516 22008 22568
rect 22060 22516 22066 22568
rect 22186 22516 22192 22568
rect 22244 22516 22250 22568
rect 20714 22488 20720 22500
rect 18693 22451 18751 22457
rect 19306 22460 20720 22488
rect 19306 22420 19334 22460
rect 20714 22448 20720 22460
rect 20772 22448 20778 22500
rect 17828 22392 19334 22420
rect 17828 22380 17834 22392
rect 19886 22380 19892 22432
rect 19944 22420 19950 22432
rect 21082 22420 21088 22432
rect 19944 22392 21088 22420
rect 19944 22380 19950 22392
rect 21082 22380 21088 22392
rect 21140 22380 21146 22432
rect 22094 22380 22100 22432
rect 22152 22380 22158 22432
rect 552 22330 23368 22352
rect 552 22278 19022 22330
rect 19074 22278 19086 22330
rect 19138 22278 19150 22330
rect 19202 22278 19214 22330
rect 19266 22278 19278 22330
rect 19330 22278 23368 22330
rect 552 22256 23368 22278
rect 4890 22176 4896 22228
rect 4948 22176 4954 22228
rect 8018 22216 8024 22228
rect 6564 22188 8024 22216
rect 4338 22108 4344 22160
rect 4396 22148 4402 22160
rect 4908 22148 4936 22176
rect 5905 22151 5963 22157
rect 5905 22148 5917 22151
rect 4396 22120 4844 22148
rect 4908 22120 5917 22148
rect 4396 22108 4402 22120
rect 4816 22080 4844 22120
rect 5905 22117 5917 22120
rect 5951 22117 5963 22151
rect 5905 22111 5963 22117
rect 6273 22151 6331 22157
rect 6273 22117 6285 22151
rect 6319 22148 6331 22151
rect 6564 22148 6592 22188
rect 8018 22176 8024 22188
rect 8076 22176 8082 22228
rect 9030 22176 9036 22228
rect 9088 22216 9094 22228
rect 9950 22216 9956 22228
rect 9088 22188 9956 22216
rect 9088 22176 9094 22188
rect 9950 22176 9956 22188
rect 10008 22176 10014 22228
rect 10137 22219 10195 22225
rect 10137 22185 10149 22219
rect 10183 22216 10195 22219
rect 10502 22216 10508 22228
rect 10183 22188 10508 22216
rect 10183 22185 10195 22188
rect 10137 22179 10195 22185
rect 10502 22176 10508 22188
rect 10560 22176 10566 22228
rect 11517 22219 11575 22225
rect 10888 22188 11468 22216
rect 6730 22148 6736 22160
rect 6319 22120 6592 22148
rect 6691 22120 6736 22148
rect 6319 22117 6331 22120
rect 6273 22111 6331 22117
rect 6730 22108 6736 22120
rect 6788 22108 6794 22160
rect 7466 22108 7472 22160
rect 7524 22148 7530 22160
rect 7524 22120 7630 22148
rect 7524 22108 7530 22120
rect 5261 22083 5319 22089
rect 5261 22080 5273 22083
rect 4816 22052 5273 22080
rect 5261 22049 5273 22052
rect 5307 22049 5319 22083
rect 5261 22043 5319 22049
rect 6089 22083 6147 22089
rect 6089 22049 6101 22083
rect 6135 22080 6147 22083
rect 6641 22083 6699 22089
rect 6135 22052 6500 22080
rect 6135 22049 6147 22052
rect 6089 22043 6147 22049
rect 6472 22024 6500 22052
rect 6641 22049 6653 22083
rect 6687 22049 6699 22083
rect 6748 22080 6776 22108
rect 7602 22089 7630 22120
rect 7834 22108 7840 22160
rect 7892 22148 7898 22160
rect 10888 22148 10916 22188
rect 11057 22151 11115 22157
rect 11057 22148 11069 22151
rect 7892 22120 10916 22148
rect 11015 22120 11069 22148
rect 7892 22108 7898 22120
rect 11057 22117 11069 22120
rect 11103 22148 11115 22151
rect 11330 22148 11336 22160
rect 11103 22120 11336 22148
rect 11103 22117 11115 22120
rect 11057 22111 11115 22117
rect 6825 22083 6883 22089
rect 6825 22080 6837 22083
rect 6748 22052 6837 22080
rect 6641 22043 6699 22049
rect 6825 22049 6837 22052
rect 6871 22049 6883 22083
rect 6825 22043 6883 22049
rect 7009 22083 7067 22089
rect 7009 22049 7021 22083
rect 7055 22049 7067 22083
rect 7009 22043 7067 22049
rect 7101 22083 7159 22089
rect 7101 22049 7113 22083
rect 7147 22049 7159 22083
rect 7101 22043 7159 22049
rect 7193 22083 7251 22089
rect 7193 22049 7205 22083
rect 7239 22049 7251 22083
rect 7193 22043 7251 22049
rect 7561 22083 7630 22089
rect 7561 22049 7573 22083
rect 7607 22052 7630 22083
rect 7607 22049 7619 22052
rect 7561 22043 7619 22049
rect 6365 22015 6423 22021
rect 6365 21981 6377 22015
rect 6411 21981 6423 22015
rect 6365 21975 6423 21981
rect 6380 21944 6408 21975
rect 6454 21972 6460 22024
rect 6512 21972 6518 22024
rect 6656 22012 6684 22043
rect 7024 22012 7052 22043
rect 6656 21984 7052 22012
rect 6840 21956 6868 21984
rect 6380 21916 6776 21944
rect 6380 21888 6408 21916
rect 5166 21836 5172 21888
rect 5224 21876 5230 21888
rect 5353 21879 5411 21885
rect 5353 21876 5365 21879
rect 5224 21848 5365 21876
rect 5224 21836 5230 21848
rect 5353 21845 5365 21848
rect 5399 21845 5411 21879
rect 5353 21839 5411 21845
rect 6362 21836 6368 21888
rect 6420 21836 6426 21888
rect 6454 21836 6460 21888
rect 6512 21836 6518 21888
rect 6748 21876 6776 21916
rect 6822 21904 6828 21956
rect 6880 21904 6886 21956
rect 7116 21876 7144 22043
rect 7208 21888 7236 22043
rect 7742 22040 7748 22092
rect 7800 22040 7806 22092
rect 8665 22083 8723 22089
rect 8665 22049 8677 22083
rect 8711 22080 8723 22083
rect 9214 22080 9220 22092
rect 8711 22052 9220 22080
rect 8711 22049 8723 22052
rect 8665 22043 8723 22049
rect 9214 22040 9220 22052
rect 9272 22040 9278 22092
rect 9309 22083 9367 22089
rect 9309 22049 9321 22083
rect 9355 22080 9367 22083
rect 9766 22080 9772 22092
rect 9355 22052 9772 22080
rect 9355 22049 9367 22052
rect 9309 22043 9367 22049
rect 9766 22040 9772 22052
rect 9824 22040 9830 22092
rect 9861 22083 9919 22089
rect 9861 22049 9873 22083
rect 9907 22049 9919 22083
rect 9861 22043 9919 22049
rect 7469 22015 7527 22021
rect 7469 21981 7481 22015
rect 7515 22012 7527 22015
rect 8478 22012 8484 22024
rect 7515 21984 8484 22012
rect 7515 21981 7527 21984
rect 7469 21975 7527 21981
rect 8478 21972 8484 21984
rect 8536 21972 8542 22024
rect 9876 22012 9904 22043
rect 9950 22040 9956 22092
rect 10008 22040 10014 22092
rect 10229 22083 10287 22089
rect 10229 22080 10241 22083
rect 10060 22052 10241 22080
rect 10060 22012 10088 22052
rect 10229 22049 10241 22052
rect 10275 22049 10287 22083
rect 10229 22043 10287 22049
rect 9692 21984 10088 22012
rect 7282 21904 7288 21956
rect 7340 21944 7346 21956
rect 7834 21944 7840 21956
rect 7340 21916 7840 21944
rect 7340 21904 7346 21916
rect 7834 21904 7840 21916
rect 7892 21904 7898 21956
rect 8496 21944 8524 21972
rect 9692 21944 9720 21984
rect 10134 21972 10140 22024
rect 10192 21972 10198 22024
rect 10689 22015 10747 22021
rect 10689 21981 10701 22015
rect 10735 22012 10747 22015
rect 11072 22012 11100 22111
rect 11330 22108 11336 22120
rect 11388 22108 11394 22160
rect 11440 22148 11468 22188
rect 11517 22185 11529 22219
rect 11563 22216 11575 22219
rect 11974 22216 11980 22228
rect 11563 22188 11980 22216
rect 11563 22185 11575 22188
rect 11517 22179 11575 22185
rect 11974 22176 11980 22188
rect 12032 22176 12038 22228
rect 12636 22188 14780 22216
rect 12636 22148 12664 22188
rect 11440 22120 12664 22148
rect 12713 22151 12771 22157
rect 12713 22117 12725 22151
rect 12759 22148 12771 22151
rect 12759 22120 12848 22148
rect 12759 22117 12771 22120
rect 12713 22111 12771 22117
rect 11514 22040 11520 22092
rect 11572 22080 11578 22092
rect 11698 22080 11704 22092
rect 11572 22052 11704 22080
rect 11572 22040 11578 22052
rect 11698 22040 11704 22052
rect 11756 22040 11762 22092
rect 12069 22083 12127 22089
rect 12069 22049 12081 22083
rect 12115 22080 12127 22083
rect 12820 22080 12848 22120
rect 13078 22108 13084 22160
rect 13136 22108 13142 22160
rect 14752 22148 14780 22188
rect 17862 22176 17868 22228
rect 17920 22216 17926 22228
rect 18598 22216 18604 22228
rect 17920 22188 18604 22216
rect 17920 22176 17926 22188
rect 18598 22176 18604 22188
rect 18656 22176 18662 22228
rect 20990 22216 20996 22228
rect 20548 22188 20996 22216
rect 15016 22160 15068 22166
rect 20548 22160 20576 22188
rect 20990 22176 20996 22188
rect 21048 22176 21054 22228
rect 21913 22219 21971 22225
rect 21913 22185 21925 22219
rect 21959 22216 21971 22219
rect 22002 22216 22008 22228
rect 21959 22188 22008 22216
rect 21959 22185 21971 22188
rect 21913 22179 21971 22185
rect 14752 22120 15016 22148
rect 17586 22108 17592 22160
rect 17644 22148 17650 22160
rect 17773 22151 17831 22157
rect 17773 22148 17785 22151
rect 17644 22120 17785 22148
rect 17644 22108 17650 22120
rect 17773 22117 17785 22120
rect 17819 22117 17831 22151
rect 18509 22151 18567 22157
rect 17773 22111 17831 22117
rect 17880 22120 18368 22148
rect 15016 22102 15068 22108
rect 12115 22052 12434 22080
rect 12820 22052 12940 22080
rect 12115 22049 12127 22052
rect 12069 22043 12127 22049
rect 10735 21984 11100 22012
rect 10735 21981 10747 21984
rect 10689 21975 10747 21981
rect 8496 21916 9720 21944
rect 10502 21904 10508 21956
rect 10560 21904 10566 21956
rect 11422 21904 11428 21956
rect 11480 21904 11486 21956
rect 6748 21848 7144 21876
rect 7190 21836 7196 21888
rect 7248 21836 7254 21888
rect 7653 21879 7711 21885
rect 7653 21845 7665 21879
rect 7699 21876 7711 21879
rect 8110 21876 8116 21888
rect 7699 21848 8116 21876
rect 7699 21845 7711 21848
rect 7653 21839 7711 21845
rect 8110 21836 8116 21848
rect 8168 21836 8174 21888
rect 8202 21836 8208 21888
rect 8260 21836 8266 21888
rect 12406 21876 12434 22052
rect 12912 22012 12940 22052
rect 13556 22012 13584 22066
rect 14458 22040 14464 22092
rect 14516 22040 14522 22092
rect 14642 22040 14648 22092
rect 14700 22080 14706 22092
rect 14737 22083 14795 22089
rect 14737 22080 14749 22083
rect 14700 22052 14749 22080
rect 14700 22040 14706 22052
rect 14737 22049 14749 22052
rect 14783 22049 14795 22083
rect 14737 22043 14795 22049
rect 16114 22040 16120 22092
rect 16172 22040 16178 22092
rect 16945 22083 17003 22089
rect 16945 22049 16957 22083
rect 16991 22080 17003 22083
rect 17034 22080 17040 22092
rect 16991 22052 17040 22080
rect 16991 22049 17003 22052
rect 16945 22043 17003 22049
rect 17034 22040 17040 22052
rect 17092 22040 17098 22092
rect 17494 22040 17500 22092
rect 17552 22040 17558 22092
rect 17681 22083 17739 22089
rect 17681 22049 17693 22083
rect 17727 22080 17739 22083
rect 17880 22080 17908 22120
rect 18340 22089 18368 22120
rect 18509 22117 18521 22151
rect 18555 22148 18567 22151
rect 19610 22148 19616 22160
rect 18555 22120 19616 22148
rect 18555 22117 18567 22120
rect 18509 22111 18567 22117
rect 19610 22108 19616 22120
rect 19668 22108 19674 22160
rect 19978 22108 19984 22160
rect 20036 22108 20042 22160
rect 20530 22148 20536 22160
rect 20088 22120 20536 22148
rect 17727 22052 17908 22080
rect 17957 22083 18015 22089
rect 17727 22049 17739 22052
rect 17681 22043 17739 22049
rect 17957 22049 17969 22083
rect 18003 22049 18015 22083
rect 18233 22083 18291 22089
rect 18233 22080 18245 22083
rect 17957 22043 18015 22049
rect 18156 22052 18245 22080
rect 12912 21984 13584 22012
rect 13556 21944 13584 21984
rect 13633 22015 13691 22021
rect 13633 21981 13645 22015
rect 13679 22012 13691 22015
rect 14274 22012 14280 22024
rect 13679 21984 14280 22012
rect 13679 21981 13691 21984
rect 13633 21975 13691 21981
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 16853 22015 16911 22021
rect 16853 21981 16865 22015
rect 16899 22012 16911 22015
rect 17696 22012 17724 22043
rect 16899 21984 16988 22012
rect 16899 21981 16911 21984
rect 16853 21975 16911 21981
rect 13556 21916 14780 21944
rect 14752 21888 14780 21916
rect 16960 21888 16988 21984
rect 17144 21984 17724 22012
rect 17144 21888 17172 21984
rect 17862 21972 17868 22024
rect 17920 22012 17926 22024
rect 17972 22012 18000 22043
rect 17920 21984 18000 22012
rect 17920 21972 17926 21984
rect 18156 21888 18184 22052
rect 18233 22049 18245 22052
rect 18279 22049 18291 22083
rect 18233 22043 18291 22049
rect 18325 22083 18383 22089
rect 18325 22049 18337 22083
rect 18371 22080 18383 22083
rect 18601 22083 18659 22089
rect 18371 22052 18425 22080
rect 18371 22049 18383 22052
rect 18325 22043 18383 22049
rect 18601 22049 18613 22083
rect 18647 22080 18659 22083
rect 18690 22080 18696 22092
rect 18647 22052 18696 22080
rect 18647 22049 18659 22052
rect 18601 22043 18659 22049
rect 18340 22012 18368 22043
rect 18690 22040 18696 22052
rect 18748 22040 18754 22092
rect 18782 22040 18788 22092
rect 18840 22080 18846 22092
rect 19061 22083 19119 22089
rect 19061 22080 19073 22083
rect 18840 22052 19073 22080
rect 18840 22040 18846 22052
rect 19061 22049 19073 22052
rect 19107 22049 19119 22083
rect 19061 22043 19119 22049
rect 19426 22040 19432 22092
rect 19484 22040 19490 22092
rect 19518 22040 19524 22092
rect 19576 22080 19582 22092
rect 19702 22080 19708 22092
rect 19576 22052 19708 22080
rect 19576 22040 19582 22052
rect 19702 22040 19708 22052
rect 19760 22080 19766 22092
rect 20088 22080 20116 22120
rect 20530 22108 20536 22120
rect 20588 22108 20594 22160
rect 20732 22120 21680 22148
rect 19760 22052 20116 22080
rect 19760 22040 19766 22052
rect 20162 22040 20168 22092
rect 20220 22040 20226 22092
rect 20254 22040 20260 22092
rect 20312 22080 20318 22092
rect 20349 22083 20407 22089
rect 20349 22080 20361 22083
rect 20312 22052 20361 22080
rect 20312 22040 20318 22052
rect 20349 22049 20361 22052
rect 20395 22049 20407 22083
rect 20349 22043 20407 22049
rect 20441 22083 20499 22089
rect 20441 22049 20453 22083
rect 20487 22080 20499 22083
rect 20548 22080 20576 22108
rect 20732 22092 20760 22120
rect 20487 22052 20576 22080
rect 20487 22049 20499 22052
rect 20441 22043 20499 22049
rect 20714 22040 20720 22092
rect 20772 22040 20778 22092
rect 21450 22040 21456 22092
rect 21508 22040 21514 22092
rect 21652 22089 21680 22120
rect 21545 22083 21603 22089
rect 21545 22049 21557 22083
rect 21591 22049 21603 22083
rect 21545 22043 21603 22049
rect 21637 22083 21695 22089
rect 21637 22049 21649 22083
rect 21683 22080 21695 22083
rect 21928 22080 21956 22179
rect 22002 22176 22008 22188
rect 22060 22176 22066 22228
rect 22186 22176 22192 22228
rect 22244 22216 22250 22228
rect 22465 22219 22523 22225
rect 22465 22216 22477 22219
rect 22244 22188 22477 22216
rect 22244 22176 22250 22188
rect 22465 22185 22477 22188
rect 22511 22185 22523 22219
rect 22465 22179 22523 22185
rect 21683 22052 21717 22080
rect 21836 22052 21956 22080
rect 21683 22049 21695 22052
rect 21637 22043 21695 22049
rect 19334 22012 19340 22024
rect 18340 21984 19340 22012
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 19889 22015 19947 22021
rect 19889 21981 19901 22015
rect 19935 22012 19947 22015
rect 20622 22012 20628 22024
rect 19935 21984 20628 22012
rect 19935 21981 19947 21984
rect 19889 21975 19947 21981
rect 20622 21972 20628 21984
rect 20680 21972 20686 22024
rect 20806 21972 20812 22024
rect 20864 22012 20870 22024
rect 21560 22012 21588 22043
rect 20864 21984 21588 22012
rect 21729 22015 21787 22021
rect 20864 21972 20870 21984
rect 21729 21981 21741 22015
rect 21775 22012 21787 22015
rect 21836 22012 21864 22052
rect 21775 21984 21864 22012
rect 21775 21981 21787 21984
rect 21729 21975 21787 21981
rect 21910 21972 21916 22024
rect 21968 22012 21974 22024
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 21968 21984 22385 22012
rect 21968 21972 21974 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 22925 22015 22983 22021
rect 22925 21981 22937 22015
rect 22971 21981 22983 22015
rect 22925 21975 22983 21981
rect 18509 21947 18567 21953
rect 18509 21913 18521 21947
rect 18555 21944 18567 21947
rect 20254 21944 20260 21956
rect 18555 21916 20260 21944
rect 18555 21913 18567 21916
rect 18509 21907 18567 21913
rect 20254 21904 20260 21916
rect 20312 21904 20318 21956
rect 22097 21947 22155 21953
rect 22097 21944 22109 21947
rect 20456 21916 22109 21944
rect 12710 21876 12716 21888
rect 12406 21848 12716 21876
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 14734 21836 14740 21888
rect 14792 21836 14798 21888
rect 16942 21836 16948 21888
rect 17000 21836 17006 21888
rect 17126 21836 17132 21888
rect 17184 21836 17190 21888
rect 17402 21836 17408 21888
rect 17460 21836 17466 21888
rect 18138 21836 18144 21888
rect 18196 21836 18202 21888
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 20456 21876 20484 21916
rect 22097 21913 22109 21916
rect 22143 21913 22155 21947
rect 22388 21944 22416 21975
rect 22557 21947 22615 21953
rect 22557 21944 22569 21947
rect 22388 21916 22569 21944
rect 22097 21907 22155 21913
rect 22557 21913 22569 21916
rect 22603 21913 22615 21947
rect 22557 21907 22615 21913
rect 19484 21848 20484 21876
rect 19484 21836 19490 21848
rect 20714 21836 20720 21888
rect 20772 21836 20778 21888
rect 21082 21836 21088 21888
rect 21140 21876 21146 21888
rect 21269 21879 21327 21885
rect 21269 21876 21281 21879
rect 21140 21848 21281 21876
rect 21140 21836 21146 21848
rect 21269 21845 21281 21848
rect 21315 21845 21327 21879
rect 22112 21876 22140 21907
rect 22940 21876 22968 21975
rect 22112 21848 22968 21876
rect 21269 21839 21327 21845
rect 552 21786 23368 21808
rect 552 21734 3662 21786
rect 3714 21734 3726 21786
rect 3778 21734 3790 21786
rect 3842 21734 3854 21786
rect 3906 21734 3918 21786
rect 3970 21734 23368 21786
rect 552 21712 23368 21734
rect 6822 21632 6828 21684
rect 6880 21632 6886 21684
rect 7282 21632 7288 21684
rect 7340 21632 7346 21684
rect 7742 21672 7748 21684
rect 7392 21644 7748 21672
rect 7300 21536 7328 21632
rect 7024 21508 7328 21536
rect 7024 21477 7052 21508
rect 7392 21480 7420 21644
rect 7742 21632 7748 21644
rect 7800 21632 7806 21684
rect 8205 21675 8263 21681
rect 8205 21641 8217 21675
rect 8251 21672 8263 21675
rect 9674 21672 9680 21684
rect 8251 21644 9680 21672
rect 8251 21641 8263 21644
rect 8205 21635 8263 21641
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 10152 21644 10824 21672
rect 7650 21564 7656 21616
rect 7708 21564 7714 21616
rect 7926 21564 7932 21616
rect 7984 21604 7990 21616
rect 8113 21607 8171 21613
rect 8113 21604 8125 21607
rect 7984 21576 8125 21604
rect 7984 21564 7990 21576
rect 8113 21573 8125 21576
rect 8159 21573 8171 21607
rect 10042 21604 10048 21616
rect 8113 21567 8171 21573
rect 8772 21576 10048 21604
rect 7009 21471 7067 21477
rect 7009 21437 7021 21471
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 7190 21428 7196 21480
rect 7248 21428 7254 21480
rect 7285 21471 7343 21477
rect 7285 21437 7297 21471
rect 7331 21468 7343 21471
rect 7374 21468 7380 21480
rect 7331 21440 7380 21468
rect 7331 21437 7343 21440
rect 7285 21431 7343 21437
rect 7374 21428 7380 21440
rect 7432 21428 7438 21480
rect 7469 21471 7527 21477
rect 7469 21437 7481 21471
rect 7515 21468 7527 21471
rect 7668 21468 7696 21564
rect 7742 21496 7748 21548
rect 7800 21536 7806 21548
rect 7837 21539 7895 21545
rect 7837 21536 7849 21539
rect 7800 21508 7849 21536
rect 7800 21496 7806 21508
rect 7837 21505 7849 21508
rect 7883 21536 7895 21539
rect 8772 21536 8800 21576
rect 10042 21564 10048 21576
rect 10100 21564 10106 21616
rect 7883 21508 8800 21536
rect 7883 21505 7895 21508
rect 7837 21499 7895 21505
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 7515 21440 7941 21468
rect 7515 21437 7527 21440
rect 7469 21431 7527 21437
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 8205 21471 8263 21477
rect 8205 21468 8217 21471
rect 7929 21431 7987 21437
rect 8036 21440 8217 21468
rect 6822 21360 6828 21412
rect 6880 21400 6886 21412
rect 7208 21400 7236 21428
rect 8036 21412 8064 21440
rect 8205 21437 8217 21440
rect 8251 21437 8263 21471
rect 8205 21431 8263 21437
rect 9490 21428 9496 21480
rect 9548 21468 9554 21480
rect 9585 21471 9643 21477
rect 9585 21468 9597 21471
rect 9548 21440 9597 21468
rect 9548 21428 9554 21440
rect 9585 21437 9597 21440
rect 9631 21468 9643 21471
rect 10152 21468 10180 21644
rect 10226 21564 10232 21616
rect 10284 21604 10290 21616
rect 10689 21607 10747 21613
rect 10689 21604 10701 21607
rect 10284 21576 10701 21604
rect 10284 21564 10290 21576
rect 10689 21573 10701 21576
rect 10735 21573 10747 21607
rect 10796 21604 10824 21644
rect 13906 21632 13912 21684
rect 13964 21632 13970 21684
rect 17126 21632 17132 21684
rect 17184 21632 17190 21684
rect 19426 21672 19432 21684
rect 17236 21644 19432 21672
rect 10796 21576 13676 21604
rect 10689 21567 10747 21573
rect 10244 21508 12388 21536
rect 10244 21477 10272 21508
rect 9631 21440 10180 21468
rect 10229 21471 10287 21477
rect 9631 21437 9643 21440
rect 9585 21431 9643 21437
rect 10229 21437 10241 21471
rect 10275 21437 10287 21471
rect 10229 21431 10287 21437
rect 8760 21412 8812 21418
rect 7653 21403 7711 21409
rect 7653 21400 7665 21403
rect 6880 21372 7665 21400
rect 6880 21360 6886 21372
rect 7653 21369 7665 21372
rect 7699 21369 7711 21403
rect 7653 21363 7711 21369
rect 8018 21360 8024 21412
rect 8076 21360 8082 21412
rect 9766 21360 9772 21412
rect 9824 21400 9830 21412
rect 10244 21400 10272 21431
rect 11146 21428 11152 21480
rect 11204 21428 11210 21480
rect 12360 21468 12388 21508
rect 12434 21496 12440 21548
rect 12492 21496 12498 21548
rect 12526 21496 12532 21548
rect 12584 21536 12590 21548
rect 13648 21536 13676 21576
rect 13924 21536 13952 21632
rect 14274 21564 14280 21616
rect 14332 21604 14338 21616
rect 16942 21604 16948 21616
rect 14332 21576 16948 21604
rect 14332 21564 14338 21576
rect 12584 21508 12756 21536
rect 12584 21496 12590 21508
rect 12728 21477 12756 21508
rect 13648 21508 13952 21536
rect 12713 21471 12771 21477
rect 9824 21372 10272 21400
rect 9824 21360 9830 21372
rect 10410 21360 10416 21412
rect 10468 21360 10474 21412
rect 10962 21360 10968 21412
rect 11020 21400 11026 21412
rect 11256 21400 11284 21454
rect 12360 21440 12572 21468
rect 11020 21372 11284 21400
rect 12161 21403 12219 21409
rect 11020 21360 11026 21372
rect 12161 21369 12173 21403
rect 12207 21400 12219 21403
rect 12544 21400 12572 21440
rect 12713 21437 12725 21471
rect 12759 21437 12771 21471
rect 13648 21470 13676 21508
rect 12713 21431 12771 21437
rect 13556 21442 13676 21470
rect 13556 21409 13584 21442
rect 13814 21428 13820 21480
rect 13872 21428 13878 21480
rect 13906 21428 13912 21480
rect 13964 21468 13970 21480
rect 14568 21477 14596 21576
rect 16942 21564 16948 21576
rect 17000 21604 17006 21616
rect 17236 21604 17264 21644
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 19521 21675 19579 21681
rect 19521 21641 19533 21675
rect 19567 21641 19579 21675
rect 19521 21635 19579 21641
rect 19705 21675 19763 21681
rect 19705 21641 19717 21675
rect 19751 21672 19763 21675
rect 20162 21672 20168 21684
rect 19751 21644 20168 21672
rect 19751 21641 19763 21644
rect 19705 21635 19763 21641
rect 17770 21604 17776 21616
rect 17000 21576 17264 21604
rect 17328 21576 17776 21604
rect 17000 21564 17006 21576
rect 14734 21496 14740 21548
rect 14792 21496 14798 21548
rect 17328 21536 17356 21576
rect 17770 21564 17776 21576
rect 17828 21564 17834 21616
rect 18138 21604 18144 21616
rect 18064 21576 18144 21604
rect 16408 21508 17356 21536
rect 17681 21539 17739 21545
rect 14185 21471 14243 21477
rect 14185 21468 14197 21471
rect 13964 21440 14197 21468
rect 13964 21428 13970 21440
rect 14185 21437 14197 21440
rect 14231 21437 14243 21471
rect 14185 21431 14243 21437
rect 14553 21471 14611 21477
rect 14553 21437 14565 21471
rect 14599 21437 14611 21471
rect 14553 21431 14611 21437
rect 15473 21471 15531 21477
rect 15473 21437 15485 21471
rect 15519 21437 15531 21471
rect 15473 21431 15531 21437
rect 13541 21403 13599 21409
rect 12207 21372 12434 21400
rect 12544 21372 13492 21400
rect 12207 21369 12219 21372
rect 12161 21363 12219 21369
rect 8760 21354 8812 21360
rect 6178 21292 6184 21344
rect 6236 21332 6242 21344
rect 7193 21335 7251 21341
rect 7193 21332 7205 21335
rect 6236 21304 7205 21332
rect 6236 21292 6242 21304
rect 7193 21301 7205 21304
rect 7239 21332 7251 21335
rect 7466 21332 7472 21344
rect 7239 21304 7472 21332
rect 7239 21301 7251 21304
rect 7193 21295 7251 21301
rect 7466 21292 7472 21304
rect 7524 21292 7530 21344
rect 10870 21292 10876 21344
rect 10928 21292 10934 21344
rect 12406 21332 12434 21372
rect 12710 21332 12716 21344
rect 12406 21304 12716 21332
rect 12710 21292 12716 21304
rect 12768 21292 12774 21344
rect 13262 21292 13268 21344
rect 13320 21332 13326 21344
rect 13357 21335 13415 21341
rect 13357 21332 13369 21335
rect 13320 21304 13369 21332
rect 13320 21292 13326 21304
rect 13357 21301 13369 21304
rect 13403 21301 13415 21335
rect 13464 21332 13492 21372
rect 13541 21369 13553 21403
rect 13587 21369 13599 21403
rect 13541 21363 13599 21369
rect 13998 21360 14004 21412
rect 14056 21360 14062 21412
rect 14642 21400 14648 21412
rect 14200 21372 14648 21400
rect 13633 21335 13691 21341
rect 13633 21332 13645 21335
rect 13464 21304 13645 21332
rect 13357 21295 13415 21301
rect 13633 21301 13645 21304
rect 13679 21332 13691 21335
rect 14200 21332 14228 21372
rect 14642 21360 14648 21372
rect 14700 21400 14706 21412
rect 15488 21400 15516 21431
rect 15562 21428 15568 21480
rect 15620 21468 15626 21480
rect 16209 21471 16267 21477
rect 16209 21468 16221 21471
rect 15620 21440 16221 21468
rect 15620 21428 15626 21440
rect 16209 21437 16221 21440
rect 16255 21468 16267 21471
rect 16408 21468 16436 21508
rect 17681 21505 17693 21539
rect 17727 21536 17739 21539
rect 17865 21539 17923 21545
rect 17865 21536 17877 21539
rect 17727 21508 17877 21536
rect 17727 21505 17739 21508
rect 17681 21499 17739 21505
rect 17865 21505 17877 21508
rect 17911 21505 17923 21539
rect 17865 21499 17923 21505
rect 16255 21440 16436 21468
rect 16255 21437 16267 21440
rect 16209 21431 16267 21437
rect 16574 21428 16580 21480
rect 16632 21468 16638 21480
rect 16853 21471 16911 21477
rect 16853 21468 16865 21471
rect 16632 21440 16865 21468
rect 16632 21428 16638 21440
rect 16853 21437 16865 21440
rect 16899 21437 16911 21471
rect 17129 21471 17187 21477
rect 17129 21468 17141 21471
rect 16853 21431 16911 21437
rect 16960 21440 17141 21468
rect 14700 21372 15516 21400
rect 15764 21372 15870 21400
rect 14700 21360 14706 21372
rect 15764 21344 15792 21372
rect 16482 21360 16488 21412
rect 16540 21400 16546 21412
rect 16960 21400 16988 21440
rect 17129 21437 17141 21440
rect 17175 21437 17187 21471
rect 17129 21431 17187 21437
rect 17586 21428 17592 21480
rect 17644 21428 17650 21480
rect 18064 21477 18092 21576
rect 18138 21564 18144 21576
rect 18196 21604 18202 21616
rect 19536 21604 19564 21635
rect 20162 21632 20168 21644
rect 20220 21632 20226 21684
rect 20901 21675 20959 21681
rect 20901 21641 20913 21675
rect 20947 21672 20959 21675
rect 20990 21672 20996 21684
rect 20947 21644 20996 21672
rect 20947 21641 20959 21644
rect 20901 21635 20959 21641
rect 20990 21632 20996 21644
rect 21048 21632 21054 21684
rect 21085 21675 21143 21681
rect 21085 21641 21097 21675
rect 21131 21672 21143 21675
rect 21266 21672 21272 21684
rect 21131 21644 21272 21672
rect 21131 21641 21143 21644
rect 21085 21635 21143 21641
rect 21266 21632 21272 21644
rect 21324 21632 21330 21684
rect 18196 21576 19564 21604
rect 18196 21564 18202 21576
rect 19978 21564 19984 21616
rect 20036 21564 20042 21616
rect 20073 21607 20131 21613
rect 20073 21573 20085 21607
rect 20119 21573 20131 21607
rect 21913 21607 21971 21613
rect 20073 21567 20131 21573
rect 20548 21576 21496 21604
rect 18690 21496 18696 21548
rect 18748 21496 18754 21548
rect 19153 21539 19211 21545
rect 19153 21505 19165 21539
rect 19199 21536 19211 21539
rect 19996 21536 20024 21564
rect 19199 21508 20024 21536
rect 19199 21505 19211 21508
rect 19153 21499 19211 21505
rect 17773 21471 17831 21477
rect 17773 21437 17785 21471
rect 17819 21468 17831 21471
rect 18049 21471 18107 21477
rect 17819 21440 17908 21468
rect 17819 21437 17831 21440
rect 17773 21431 17831 21437
rect 17880 21412 17908 21440
rect 18049 21437 18061 21471
rect 18095 21437 18107 21471
rect 18049 21431 18107 21437
rect 18782 21428 18788 21480
rect 18840 21468 18846 21480
rect 19061 21471 19119 21477
rect 19061 21468 19073 21471
rect 18840 21440 19073 21468
rect 18840 21428 18846 21440
rect 19061 21437 19073 21440
rect 19107 21468 19119 21471
rect 19107 21440 19748 21468
rect 19107 21437 19119 21440
rect 19061 21431 19119 21437
rect 16540 21372 16988 21400
rect 17037 21403 17095 21409
rect 16540 21360 16546 21372
rect 17037 21369 17049 21403
rect 17083 21369 17095 21403
rect 17037 21363 17095 21369
rect 13679 21304 14228 21332
rect 13679 21301 13691 21304
rect 13633 21295 13691 21301
rect 14274 21292 14280 21344
rect 14332 21292 14338 21344
rect 14918 21292 14924 21344
rect 14976 21332 14982 21344
rect 15746 21332 15752 21344
rect 14976 21304 15752 21332
rect 14976 21292 14982 21304
rect 15746 21292 15752 21304
rect 15804 21292 15810 21344
rect 16666 21292 16672 21344
rect 16724 21332 16730 21344
rect 17052 21332 17080 21363
rect 17862 21360 17868 21412
rect 17920 21360 17926 21412
rect 19334 21360 19340 21412
rect 19392 21360 19398 21412
rect 19518 21360 19524 21412
rect 19576 21409 19582 21412
rect 19576 21403 19611 21409
rect 19599 21369 19611 21403
rect 19720 21400 19748 21440
rect 19794 21428 19800 21480
rect 19852 21428 19858 21480
rect 20088 21468 20116 21567
rect 20548 21548 20576 21576
rect 20530 21496 20536 21548
rect 20588 21496 20594 21548
rect 20898 21496 20904 21548
rect 20956 21536 20962 21548
rect 20956 21508 21404 21536
rect 20956 21496 20962 21508
rect 20088 21440 20944 21468
rect 19889 21403 19947 21409
rect 19889 21400 19901 21403
rect 19720 21372 19901 21400
rect 19576 21363 19611 21369
rect 19889 21369 19901 21372
rect 19935 21369 19947 21403
rect 19889 21363 19947 21369
rect 20073 21403 20131 21409
rect 20073 21369 20085 21403
rect 20119 21400 20131 21403
rect 20254 21400 20260 21412
rect 20119 21372 20260 21400
rect 20119 21369 20131 21372
rect 20073 21363 20131 21369
rect 19576 21360 19582 21363
rect 20254 21360 20260 21372
rect 20312 21360 20318 21412
rect 20530 21360 20536 21412
rect 20588 21360 20594 21412
rect 20717 21403 20775 21409
rect 20717 21369 20729 21403
rect 20763 21400 20775 21403
rect 20806 21400 20812 21412
rect 20763 21372 20812 21400
rect 20763 21369 20775 21372
rect 20717 21363 20775 21369
rect 20806 21360 20812 21372
rect 20864 21360 20870 21412
rect 20916 21400 20944 21440
rect 20990 21428 20996 21480
rect 21048 21468 21054 21480
rect 21376 21477 21404 21508
rect 21468 21477 21496 21576
rect 21913 21573 21925 21607
rect 21959 21604 21971 21607
rect 22373 21607 22431 21613
rect 21959 21576 22094 21604
rect 21959 21573 21971 21576
rect 21913 21567 21971 21573
rect 22066 21548 22094 21576
rect 22373 21573 22385 21607
rect 22419 21573 22431 21607
rect 22373 21567 22431 21573
rect 22066 21508 22100 21548
rect 22094 21496 22100 21508
rect 22152 21496 22158 21548
rect 21177 21471 21235 21477
rect 21177 21468 21189 21471
rect 21048 21440 21189 21468
rect 21048 21428 21054 21440
rect 21177 21437 21189 21440
rect 21223 21437 21235 21471
rect 21177 21431 21235 21437
rect 21361 21471 21419 21477
rect 21361 21437 21373 21471
rect 21407 21437 21419 21471
rect 21361 21431 21419 21437
rect 21453 21471 21511 21477
rect 21453 21437 21465 21471
rect 21499 21437 21511 21471
rect 22388 21468 22416 21567
rect 21453 21431 21511 21437
rect 22066 21440 22416 21468
rect 21545 21403 21603 21409
rect 21545 21400 21557 21403
rect 20916 21372 21557 21400
rect 21545 21369 21557 21372
rect 21591 21400 21603 21403
rect 22066 21400 22094 21440
rect 21591 21372 22094 21400
rect 21591 21369 21603 21372
rect 21545 21363 21603 21369
rect 16724 21304 17080 21332
rect 16724 21292 16730 21304
rect 18230 21292 18236 21344
rect 18288 21292 18294 21344
rect 20548 21332 20576 21360
rect 20917 21335 20975 21341
rect 20917 21332 20929 21335
rect 20548 21304 20929 21332
rect 20917 21301 20929 21304
rect 20963 21301 20975 21335
rect 20917 21295 20975 21301
rect 21174 21292 21180 21344
rect 21232 21332 21238 21344
rect 21275 21335 21333 21341
rect 21275 21332 21287 21335
rect 21232 21304 21287 21332
rect 21232 21292 21238 21304
rect 21275 21301 21287 21304
rect 21321 21301 21333 21335
rect 21275 21295 21333 21301
rect 22002 21292 22008 21344
rect 22060 21292 22066 21344
rect 22554 21292 22560 21344
rect 22612 21292 22618 21344
rect 552 21242 23368 21264
rect 552 21190 19022 21242
rect 19074 21190 19086 21242
rect 19138 21190 19150 21242
rect 19202 21190 19214 21242
rect 19266 21190 19278 21242
rect 19330 21190 23368 21242
rect 552 21168 23368 21190
rect 6362 21088 6368 21140
rect 6420 21128 6426 21140
rect 6457 21131 6515 21137
rect 6457 21128 6469 21131
rect 6420 21100 6469 21128
rect 6420 21088 6426 21100
rect 6457 21097 6469 21100
rect 6503 21097 6515 21131
rect 6457 21091 6515 21097
rect 7282 21088 7288 21140
rect 7340 21088 7346 21140
rect 7374 21088 7380 21140
rect 7432 21128 7438 21140
rect 8202 21128 8208 21140
rect 7432 21100 7972 21128
rect 7432 21088 7438 21100
rect 5350 21060 5356 21072
rect 4448 21032 5356 21060
rect 4341 20995 4399 21001
rect 4341 20961 4353 20995
rect 4387 20961 4399 20995
rect 4341 20955 4399 20961
rect 4356 20788 4384 20955
rect 4448 20936 4476 21032
rect 5350 21020 5356 21032
rect 5408 21020 5414 21072
rect 5552 21032 6224 21060
rect 4614 20952 4620 21004
rect 4672 20992 4678 21004
rect 5445 20995 5503 21001
rect 5445 20992 5457 20995
rect 4672 20964 5457 20992
rect 4672 20952 4678 20964
rect 5445 20961 5457 20964
rect 5491 20992 5503 20995
rect 5552 20992 5580 21032
rect 5491 20964 5580 20992
rect 5491 20961 5503 20964
rect 5445 20955 5503 20961
rect 5626 20952 5632 21004
rect 5684 20952 5690 21004
rect 5813 20995 5871 21001
rect 5813 20961 5825 20995
rect 5859 20961 5871 20995
rect 5813 20955 5871 20961
rect 4430 20884 4436 20936
rect 4488 20884 4494 20936
rect 5350 20884 5356 20936
rect 5408 20924 5414 20936
rect 5828 20924 5856 20955
rect 5994 20952 6000 21004
rect 6052 20952 6058 21004
rect 6196 21001 6224 21032
rect 6089 20995 6147 21001
rect 6089 20961 6101 20995
rect 6135 20961 6147 20995
rect 6089 20955 6147 20961
rect 6181 20995 6239 21001
rect 6181 20961 6193 20995
rect 6227 20992 6239 20995
rect 6270 20992 6276 21004
rect 6227 20964 6276 20992
rect 6227 20961 6239 20964
rect 6181 20955 6239 20961
rect 5408 20896 5856 20924
rect 5408 20884 5414 20896
rect 4709 20859 4767 20865
rect 4709 20825 4721 20859
rect 4755 20856 4767 20859
rect 5258 20856 5264 20868
rect 4755 20828 5264 20856
rect 4755 20825 4767 20828
rect 4709 20819 4767 20825
rect 5258 20816 5264 20828
rect 5316 20856 5322 20868
rect 6104 20856 6132 20955
rect 6270 20952 6276 20964
rect 6328 20952 6334 21004
rect 6362 20952 6368 21004
rect 6420 20952 6426 21004
rect 7300 21001 7328 21088
rect 7944 21004 7972 21100
rect 8036 21100 8208 21128
rect 7285 20995 7343 21001
rect 7285 20961 7297 20995
rect 7331 20961 7343 20995
rect 7285 20955 7343 20961
rect 7377 20995 7435 21001
rect 7377 20961 7389 20995
rect 7423 20992 7435 20995
rect 7466 20992 7472 21004
rect 7423 20964 7472 20992
rect 7423 20961 7435 20964
rect 7377 20955 7435 20961
rect 7466 20952 7472 20964
rect 7524 20952 7530 21004
rect 7561 20995 7619 21001
rect 7561 20961 7573 20995
rect 7607 20961 7619 20995
rect 7561 20955 7619 20961
rect 6380 20924 6408 20952
rect 6822 20924 6828 20936
rect 6380 20896 6828 20924
rect 6822 20884 6828 20896
rect 6880 20924 6886 20936
rect 7576 20924 7604 20955
rect 7926 20952 7932 21004
rect 7984 20952 7990 21004
rect 6880 20896 7604 20924
rect 6880 20884 6886 20896
rect 7650 20884 7656 20936
rect 7708 20924 7714 20936
rect 8036 20924 8064 21100
rect 8202 21088 8208 21100
rect 8260 21088 8266 21140
rect 10410 21088 10416 21140
rect 10468 21088 10474 21140
rect 10870 21088 10876 21140
rect 10928 21088 10934 21140
rect 11057 21131 11115 21137
rect 11057 21097 11069 21131
rect 11103 21128 11115 21131
rect 11146 21128 11152 21140
rect 11103 21100 11152 21128
rect 11103 21097 11115 21100
rect 11057 21091 11115 21097
rect 11146 21088 11152 21100
rect 11204 21128 11210 21140
rect 12897 21131 12955 21137
rect 11204 21100 11560 21128
rect 11204 21088 11210 21100
rect 9309 21063 9367 21069
rect 9309 21029 9321 21063
rect 9355 21060 9367 21063
rect 10428 21060 10456 21088
rect 9355 21032 10456 21060
rect 10888 21060 10916 21088
rect 10888 21032 11284 21060
rect 9355 21029 9367 21032
rect 9309 21023 9367 21029
rect 8110 20952 8116 21004
rect 8168 20992 8174 21004
rect 8481 20995 8539 21001
rect 8481 20992 8493 20995
rect 8168 20964 8493 20992
rect 8168 20952 8174 20964
rect 8481 20961 8493 20964
rect 8527 20961 8539 20995
rect 8481 20955 8539 20961
rect 10045 20995 10103 21001
rect 10045 20961 10057 20995
rect 10091 20992 10103 20995
rect 10226 20992 10232 21004
rect 10091 20964 10232 20992
rect 10091 20961 10103 20964
rect 10045 20955 10103 20961
rect 10226 20952 10232 20964
rect 10284 20952 10290 21004
rect 10321 20995 10379 21001
rect 10321 20961 10333 20995
rect 10367 20992 10379 20995
rect 10428 20992 10456 21032
rect 10367 20964 10456 20992
rect 10689 20995 10747 21001
rect 10367 20961 10379 20964
rect 10321 20955 10379 20961
rect 10689 20961 10701 20995
rect 10735 20992 10747 20995
rect 10962 20992 10968 21004
rect 10735 20964 10968 20992
rect 10735 20961 10747 20964
rect 10689 20955 10747 20961
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 11256 21001 11284 21032
rect 11241 20995 11299 21001
rect 11241 20961 11253 20995
rect 11287 20961 11299 20995
rect 11532 20992 11560 21100
rect 12897 21097 12909 21131
rect 12943 21128 12955 21131
rect 13906 21128 13912 21140
rect 12943 21100 13912 21128
rect 12943 21097 12955 21100
rect 12897 21091 12955 21097
rect 13906 21088 13912 21100
rect 13964 21088 13970 21140
rect 16298 21088 16304 21140
rect 16356 21128 16362 21140
rect 19245 21131 19303 21137
rect 16356 21100 17632 21128
rect 16356 21088 16362 21100
rect 11698 21020 11704 21072
rect 11756 21060 11762 21072
rect 13354 21069 13360 21072
rect 12437 21063 12495 21069
rect 12437 21060 12449 21063
rect 11756 21032 12449 21060
rect 11756 21020 11762 21032
rect 12437 21029 12449 21032
rect 12483 21029 12495 21063
rect 12437 21023 12495 21029
rect 13081 21063 13139 21069
rect 13081 21029 13093 21063
rect 13127 21029 13139 21063
rect 13081 21023 13139 21029
rect 13297 21063 13360 21069
rect 13297 21029 13309 21063
rect 13343 21029 13360 21063
rect 13297 21023 13360 21029
rect 12802 20992 12808 21004
rect 11532 20964 12808 20992
rect 11241 20955 11299 20961
rect 12802 20952 12808 20964
rect 12860 20952 12866 21004
rect 8389 20927 8447 20933
rect 8389 20924 8401 20927
rect 7708 20896 8401 20924
rect 7708 20884 7714 20896
rect 8389 20893 8401 20896
rect 8435 20893 8447 20927
rect 8389 20887 8447 20893
rect 11882 20884 11888 20936
rect 11940 20924 11946 20936
rect 13096 20924 13124 21023
rect 13354 21020 13360 21023
rect 13412 21020 13418 21072
rect 14642 21020 14648 21072
rect 14700 21020 14706 21072
rect 17604 21060 17632 21100
rect 19245 21097 19257 21131
rect 19291 21128 19303 21131
rect 19794 21128 19800 21140
rect 19291 21100 19800 21128
rect 19291 21097 19303 21100
rect 19245 21091 19303 21097
rect 19794 21088 19800 21100
rect 19852 21088 19858 21140
rect 19978 21088 19984 21140
rect 20036 21088 20042 21140
rect 19702 21060 19708 21072
rect 16592 21032 17540 21060
rect 17604 21032 19708 21060
rect 16592 21004 16620 21032
rect 13998 20952 14004 21004
rect 14056 20992 14062 21004
rect 14185 20995 14243 21001
rect 14185 20992 14197 20995
rect 14056 20964 14197 20992
rect 14056 20952 14062 20964
rect 14185 20961 14197 20964
rect 14231 20961 14243 20995
rect 14185 20955 14243 20961
rect 14921 20995 14979 21001
rect 14921 20961 14933 20995
rect 14967 20992 14979 20995
rect 15194 20992 15200 21004
rect 14967 20964 15200 20992
rect 14967 20961 14979 20964
rect 14921 20955 14979 20961
rect 15194 20952 15200 20964
rect 15252 20952 15258 21004
rect 15378 20952 15384 21004
rect 15436 20992 15442 21004
rect 16393 20995 16451 21001
rect 16393 20992 16405 20995
rect 15436 20964 16405 20992
rect 15436 20952 15442 20964
rect 16393 20961 16405 20964
rect 16439 20992 16451 20995
rect 16482 20992 16488 21004
rect 16439 20964 16488 20992
rect 16439 20961 16451 20964
rect 16393 20955 16451 20961
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 16574 20952 16580 21004
rect 16632 20952 16638 21004
rect 17512 21001 17540 21032
rect 19702 21020 19708 21032
rect 19760 21020 19766 21072
rect 17313 20995 17371 21001
rect 17313 20961 17325 20995
rect 17359 20961 17371 20995
rect 17313 20955 17371 20961
rect 17497 20995 17555 21001
rect 17497 20961 17509 20995
rect 17543 20992 17555 20995
rect 17586 20992 17592 21004
rect 17543 20964 17592 20992
rect 17543 20961 17555 20964
rect 17497 20955 17555 20961
rect 11940 20896 13584 20924
rect 11940 20884 11946 20896
rect 5316 20828 6132 20856
rect 7561 20859 7619 20865
rect 5316 20816 5322 20828
rect 7561 20825 7573 20859
rect 7607 20856 7619 20859
rect 8018 20856 8024 20868
rect 7607 20828 8024 20856
rect 7607 20825 7619 20828
rect 7561 20819 7619 20825
rect 8018 20816 8024 20828
rect 8076 20816 8082 20868
rect 8110 20816 8116 20868
rect 8168 20816 8174 20868
rect 12710 20816 12716 20868
rect 12768 20816 12774 20868
rect 13446 20816 13452 20868
rect 13504 20816 13510 20868
rect 13556 20856 13584 20896
rect 15746 20884 15752 20936
rect 15804 20924 15810 20936
rect 16301 20927 16359 20933
rect 16301 20924 16313 20927
rect 15804 20896 16313 20924
rect 15804 20884 15810 20896
rect 16301 20893 16313 20896
rect 16347 20924 16359 20927
rect 16666 20924 16672 20936
rect 16347 20896 16672 20924
rect 16347 20893 16359 20896
rect 16301 20887 16359 20893
rect 16666 20884 16672 20896
rect 16724 20884 16730 20936
rect 17221 20927 17279 20933
rect 17221 20893 17233 20927
rect 17267 20924 17279 20927
rect 17328 20924 17356 20955
rect 17586 20952 17592 20964
rect 17644 20952 17650 21004
rect 17954 20952 17960 21004
rect 18012 20952 18018 21004
rect 19153 20995 19211 21001
rect 19153 20961 19165 20995
rect 19199 20992 19211 20995
rect 19996 20992 20024 21088
rect 21174 21060 21180 21072
rect 20824 21032 21180 21060
rect 20824 21001 20852 21032
rect 21174 21020 21180 21032
rect 21232 21060 21238 21072
rect 21232 21032 21496 21060
rect 21232 21020 21238 21032
rect 19199 20964 20024 20992
rect 20809 20995 20867 21001
rect 19199 20961 19211 20964
rect 19153 20955 19211 20961
rect 20809 20961 20821 20995
rect 20855 20961 20867 20995
rect 20809 20955 20867 20961
rect 20993 20995 21051 21001
rect 20993 20961 21005 20995
rect 21039 20992 21051 20995
rect 21082 20992 21088 21004
rect 21039 20964 21088 20992
rect 21039 20961 21051 20964
rect 20993 20955 21051 20961
rect 21082 20952 21088 20964
rect 21140 20952 21146 21004
rect 21266 20952 21272 21004
rect 21324 20952 21330 21004
rect 21468 21001 21496 21032
rect 21453 20995 21511 21001
rect 21453 20961 21465 20995
rect 21499 20961 21511 20995
rect 21453 20955 21511 20961
rect 21729 20995 21787 21001
rect 21729 20961 21741 20995
rect 21775 20961 21787 20995
rect 21729 20955 21787 20961
rect 17972 20924 18000 20952
rect 17267 20896 18000 20924
rect 20901 20927 20959 20933
rect 17267 20893 17279 20896
rect 17221 20887 17279 20893
rect 20901 20893 20913 20927
rect 20947 20893 20959 20927
rect 21100 20924 21128 20952
rect 21744 20924 21772 20955
rect 21100 20896 21772 20924
rect 20901 20887 20959 20893
rect 14458 20856 14464 20868
rect 13556 20828 14464 20856
rect 14458 20816 14464 20828
rect 14516 20816 14522 20868
rect 17402 20816 17408 20868
rect 17460 20856 17466 20868
rect 20714 20856 20720 20868
rect 17460 20828 20720 20856
rect 17460 20816 17466 20828
rect 20714 20816 20720 20828
rect 20772 20816 20778 20868
rect 20916 20856 20944 20887
rect 21266 20856 21272 20868
rect 20916 20828 21272 20856
rect 21266 20816 21272 20828
rect 21324 20816 21330 20868
rect 5166 20788 5172 20800
rect 4356 20760 5172 20788
rect 5166 20748 5172 20760
rect 5224 20748 5230 20800
rect 5626 20748 5632 20800
rect 5684 20748 5690 20800
rect 7742 20748 7748 20800
rect 7800 20748 7806 20800
rect 11425 20791 11483 20797
rect 11425 20757 11437 20791
rect 11471 20788 11483 20791
rect 11606 20788 11612 20800
rect 11471 20760 11612 20788
rect 11471 20757 11483 20760
rect 11425 20751 11483 20757
rect 11606 20748 11612 20760
rect 11664 20748 11670 20800
rect 13265 20791 13323 20797
rect 13265 20757 13277 20791
rect 13311 20788 13323 20791
rect 14550 20788 14556 20800
rect 13311 20760 14556 20788
rect 13311 20757 13323 20760
rect 13265 20751 13323 20757
rect 14550 20748 14556 20760
rect 14608 20748 14614 20800
rect 17494 20748 17500 20800
rect 17552 20748 17558 20800
rect 20625 20791 20683 20797
rect 20625 20757 20637 20791
rect 20671 20788 20683 20791
rect 20806 20788 20812 20800
rect 20671 20760 20812 20788
rect 20671 20757 20683 20760
rect 20625 20751 20683 20757
rect 20806 20748 20812 20760
rect 20864 20748 20870 20800
rect 21910 20748 21916 20800
rect 21968 20748 21974 20800
rect 552 20698 23368 20720
rect 552 20646 3662 20698
rect 3714 20646 3726 20698
rect 3778 20646 3790 20698
rect 3842 20646 3854 20698
rect 3906 20646 3918 20698
rect 3970 20646 23368 20698
rect 552 20624 23368 20646
rect 5626 20544 5632 20596
rect 5684 20584 5690 20596
rect 5994 20584 6000 20596
rect 5684 20556 6000 20584
rect 5684 20544 5690 20556
rect 5994 20544 6000 20556
rect 6052 20544 6058 20596
rect 6365 20587 6423 20593
rect 6365 20553 6377 20587
rect 6411 20584 6423 20587
rect 7742 20584 7748 20596
rect 6411 20556 7748 20584
rect 6411 20553 6423 20556
rect 6365 20547 6423 20553
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 7926 20544 7932 20596
rect 7984 20544 7990 20596
rect 12802 20544 12808 20596
rect 12860 20584 12866 20596
rect 12897 20587 12955 20593
rect 12897 20584 12909 20587
rect 12860 20556 12909 20584
rect 12860 20544 12866 20556
rect 12897 20553 12909 20556
rect 12943 20553 12955 20587
rect 12897 20547 12955 20553
rect 15194 20544 15200 20596
rect 15252 20544 15258 20596
rect 18046 20544 18052 20596
rect 18104 20584 18110 20596
rect 18693 20587 18751 20593
rect 18693 20584 18705 20587
rect 18104 20556 18705 20584
rect 18104 20544 18110 20556
rect 18693 20553 18705 20556
rect 18739 20553 18751 20587
rect 21910 20584 21916 20596
rect 18693 20547 18751 20553
rect 21376 20556 21916 20584
rect 5077 20519 5135 20525
rect 5077 20485 5089 20519
rect 5123 20516 5135 20519
rect 5810 20516 5816 20528
rect 5123 20488 5816 20516
rect 5123 20485 5135 20488
rect 5077 20479 5135 20485
rect 5810 20476 5816 20488
rect 5868 20476 5874 20528
rect 7282 20476 7288 20528
rect 7340 20476 7346 20528
rect 4249 20451 4307 20457
rect 4249 20417 4261 20451
rect 4295 20448 4307 20451
rect 6089 20451 6147 20457
rect 6089 20448 6101 20451
rect 4295 20420 6101 20448
rect 4295 20417 4307 20420
rect 4249 20411 4307 20417
rect 6089 20417 6101 20420
rect 6135 20417 6147 20451
rect 6089 20411 6147 20417
rect 7837 20451 7895 20457
rect 7837 20417 7849 20451
rect 7883 20448 7895 20451
rect 7944 20448 7972 20544
rect 12728 20488 13492 20516
rect 7883 20420 7972 20448
rect 7883 20417 7895 20420
rect 7837 20411 7895 20417
rect 8202 20408 8208 20460
rect 8260 20408 8266 20460
rect 4157 20383 4215 20389
rect 4157 20349 4169 20383
rect 4203 20349 4215 20383
rect 4157 20343 4215 20349
rect 4172 20312 4200 20343
rect 4338 20340 4344 20392
rect 4396 20340 4402 20392
rect 4430 20340 4436 20392
rect 4488 20340 4494 20392
rect 4614 20340 4620 20392
rect 4672 20340 4678 20392
rect 4985 20383 5043 20389
rect 4985 20349 4997 20383
rect 5031 20349 5043 20383
rect 4985 20343 5043 20349
rect 4246 20312 4252 20324
rect 4172 20284 4252 20312
rect 4246 20272 4252 20284
rect 4304 20312 4310 20324
rect 4632 20312 4660 20340
rect 4304 20284 4660 20312
rect 4801 20315 4859 20321
rect 4304 20272 4310 20284
rect 4801 20281 4813 20315
rect 4847 20312 4859 20315
rect 5000 20312 5028 20343
rect 5166 20340 5172 20392
rect 5224 20340 5230 20392
rect 5258 20340 5264 20392
rect 5316 20340 5322 20392
rect 5350 20340 5356 20392
rect 5408 20340 5414 20392
rect 5537 20383 5595 20389
rect 5537 20349 5549 20383
rect 5583 20380 5595 20383
rect 5997 20383 6055 20389
rect 5997 20380 6009 20383
rect 5583 20352 6009 20380
rect 5583 20349 5595 20352
rect 5537 20343 5595 20349
rect 5997 20349 6009 20352
rect 6043 20380 6055 20383
rect 6362 20380 6368 20392
rect 6043 20352 6368 20380
rect 6043 20349 6055 20352
rect 5997 20343 6055 20349
rect 6362 20340 6368 20352
rect 6420 20340 6426 20392
rect 7650 20340 7656 20392
rect 7708 20380 7714 20392
rect 7926 20380 7932 20392
rect 7708 20352 7932 20380
rect 7708 20340 7714 20352
rect 7926 20340 7932 20352
rect 7984 20380 7990 20392
rect 8021 20383 8079 20389
rect 8021 20380 8033 20383
rect 7984 20352 8033 20380
rect 7984 20340 7990 20352
rect 8021 20349 8033 20352
rect 8067 20349 8079 20383
rect 8021 20343 8079 20349
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20380 8171 20383
rect 8220 20380 8248 20408
rect 8159 20352 8248 20380
rect 8159 20349 8171 20352
rect 8113 20343 8171 20349
rect 12158 20340 12164 20392
rect 12216 20380 12222 20392
rect 12728 20389 12756 20488
rect 13464 20460 13492 20488
rect 13173 20451 13231 20457
rect 13173 20448 13185 20451
rect 12912 20420 13185 20448
rect 12912 20389 12940 20420
rect 13173 20417 13185 20420
rect 13219 20417 13231 20451
rect 13173 20411 13231 20417
rect 13446 20408 13452 20460
rect 13504 20408 13510 20460
rect 15212 20448 15240 20544
rect 18785 20451 18843 20457
rect 18785 20448 18797 20451
rect 13740 20420 15240 20448
rect 17512 20420 18797 20448
rect 12713 20383 12771 20389
rect 12713 20380 12725 20383
rect 12216 20352 12725 20380
rect 12216 20340 12222 20352
rect 12713 20349 12725 20352
rect 12759 20349 12771 20383
rect 12713 20343 12771 20349
rect 12897 20383 12955 20389
rect 12897 20349 12909 20383
rect 12943 20349 12955 20383
rect 12897 20343 12955 20349
rect 12986 20340 12992 20392
rect 13044 20380 13050 20392
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 13044 20352 13093 20380
rect 13044 20340 13050 20352
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 13081 20343 13139 20349
rect 13265 20383 13323 20389
rect 13265 20349 13277 20383
rect 13311 20380 13323 20383
rect 13354 20380 13360 20392
rect 13311 20352 13360 20380
rect 13311 20349 13323 20352
rect 13265 20343 13323 20349
rect 4847 20284 5028 20312
rect 4847 20281 4859 20284
rect 4801 20275 4859 20281
rect 5000 20244 5028 20284
rect 5368 20244 5396 20340
rect 7009 20315 7067 20321
rect 7009 20281 7021 20315
rect 7055 20312 7067 20315
rect 7098 20312 7104 20324
rect 7055 20284 7104 20312
rect 7055 20281 7067 20284
rect 7009 20275 7067 20281
rect 7098 20272 7104 20284
rect 7156 20272 7162 20324
rect 9398 20312 9404 20324
rect 7484 20284 9404 20312
rect 5000 20216 5396 20244
rect 5718 20204 5724 20256
rect 5776 20204 5782 20256
rect 7484 20253 7512 20284
rect 9398 20272 9404 20284
rect 9456 20272 9462 20324
rect 7469 20247 7527 20253
rect 7469 20213 7481 20247
rect 7515 20213 7527 20247
rect 7469 20207 7527 20213
rect 7837 20247 7895 20253
rect 7837 20213 7849 20247
rect 7883 20244 7895 20247
rect 8386 20244 8392 20256
rect 7883 20216 8392 20244
rect 7883 20213 7895 20216
rect 7837 20207 7895 20213
rect 8386 20204 8392 20216
rect 8444 20204 8450 20256
rect 13096 20244 13124 20343
rect 13354 20340 13360 20352
rect 13412 20380 13418 20392
rect 13740 20389 13768 20420
rect 17512 20392 17540 20420
rect 18785 20417 18797 20420
rect 18831 20417 18843 20451
rect 18785 20411 18843 20417
rect 13725 20383 13783 20389
rect 13412 20352 13676 20380
rect 13412 20340 13418 20352
rect 13538 20272 13544 20324
rect 13596 20272 13602 20324
rect 13648 20312 13676 20352
rect 13725 20349 13737 20383
rect 13771 20349 13783 20383
rect 13725 20343 13783 20349
rect 13909 20383 13967 20389
rect 13909 20349 13921 20383
rect 13955 20380 13967 20383
rect 13998 20380 14004 20392
rect 13955 20352 14004 20380
rect 13955 20349 13967 20352
rect 13909 20343 13967 20349
rect 13998 20340 14004 20352
rect 14056 20340 14062 20392
rect 14369 20383 14427 20389
rect 14369 20349 14381 20383
rect 14415 20349 14427 20383
rect 14369 20343 14427 20349
rect 14384 20312 14412 20343
rect 14458 20340 14464 20392
rect 14516 20340 14522 20392
rect 14550 20340 14556 20392
rect 14608 20340 14614 20392
rect 14642 20340 14648 20392
rect 14700 20340 14706 20392
rect 14921 20383 14979 20389
rect 14921 20349 14933 20383
rect 14967 20380 14979 20383
rect 15378 20380 15384 20392
rect 14967 20352 15384 20380
rect 14967 20349 14979 20352
rect 14921 20343 14979 20349
rect 15378 20340 15384 20352
rect 15436 20380 15442 20392
rect 15749 20383 15807 20389
rect 15749 20380 15761 20383
rect 15436 20352 15761 20380
rect 15436 20340 15442 20352
rect 15749 20349 15761 20352
rect 15795 20349 15807 20383
rect 15749 20343 15807 20349
rect 16485 20383 16543 20389
rect 16485 20349 16497 20383
rect 16531 20380 16543 20383
rect 17402 20380 17408 20392
rect 16531 20352 17408 20380
rect 16531 20349 16543 20352
rect 16485 20343 16543 20349
rect 17402 20340 17408 20352
rect 17460 20340 17466 20392
rect 17494 20340 17500 20392
rect 17552 20340 17558 20392
rect 17586 20340 17592 20392
rect 17644 20340 17650 20392
rect 17954 20340 17960 20392
rect 18012 20340 18018 20392
rect 18230 20340 18236 20392
rect 18288 20380 18294 20392
rect 18693 20383 18751 20389
rect 18693 20380 18705 20383
rect 18288 20352 18705 20380
rect 18288 20340 18294 20352
rect 18693 20349 18705 20352
rect 18739 20349 18751 20383
rect 18693 20343 18751 20349
rect 20806 20340 20812 20392
rect 20864 20380 20870 20392
rect 21376 20389 21404 20556
rect 21910 20544 21916 20556
rect 21968 20544 21974 20596
rect 22002 20516 22008 20528
rect 21836 20488 22008 20516
rect 21836 20389 21864 20488
rect 22002 20476 22008 20488
rect 22060 20516 22066 20528
rect 22060 20488 22416 20516
rect 22060 20476 22066 20488
rect 21910 20408 21916 20460
rect 21968 20448 21974 20460
rect 21968 20420 22140 20448
rect 21968 20408 21974 20420
rect 22112 20389 22140 20420
rect 22388 20389 22416 20488
rect 20901 20383 20959 20389
rect 20901 20380 20913 20383
rect 20864 20352 20913 20380
rect 20864 20340 20870 20352
rect 20901 20349 20913 20352
rect 20947 20349 20959 20383
rect 20901 20343 20959 20349
rect 21085 20383 21143 20389
rect 21085 20349 21097 20383
rect 21131 20380 21143 20383
rect 21361 20383 21419 20389
rect 21361 20380 21373 20383
rect 21131 20352 21373 20380
rect 21131 20349 21143 20352
rect 21085 20343 21143 20349
rect 21361 20349 21373 20352
rect 21407 20349 21419 20383
rect 21361 20343 21419 20349
rect 21637 20383 21695 20389
rect 21637 20349 21649 20383
rect 21683 20349 21695 20383
rect 21637 20343 21695 20349
rect 21821 20383 21879 20389
rect 21821 20349 21833 20383
rect 21867 20349 21879 20383
rect 21821 20343 21879 20349
rect 22105 20383 22163 20389
rect 22105 20349 22117 20383
rect 22151 20349 22163 20383
rect 22105 20343 22163 20349
rect 22373 20383 22431 20389
rect 22373 20349 22385 20383
rect 22419 20349 22431 20383
rect 22373 20343 22431 20349
rect 14568 20312 14596 20340
rect 13648 20284 14320 20312
rect 14384 20284 14596 20312
rect 13722 20244 13728 20256
rect 13096 20216 13728 20244
rect 13722 20204 13728 20216
rect 13780 20244 13786 20256
rect 14185 20247 14243 20253
rect 14185 20244 14197 20247
rect 13780 20216 14197 20244
rect 13780 20204 13786 20216
rect 14185 20213 14197 20216
rect 14231 20213 14243 20247
rect 14292 20244 14320 20284
rect 15194 20272 15200 20324
rect 15252 20272 15258 20324
rect 20916 20312 20944 20343
rect 21652 20312 21680 20343
rect 22554 20340 22560 20392
rect 22612 20340 22618 20392
rect 21913 20315 21971 20321
rect 21913 20312 21925 20315
rect 20916 20284 21925 20312
rect 21913 20281 21925 20284
rect 21959 20281 21971 20315
rect 22465 20315 22523 20321
rect 22465 20312 22477 20315
rect 21913 20275 21971 20281
rect 22066 20284 22477 20312
rect 16298 20244 16304 20256
rect 14292 20216 16304 20244
rect 14185 20207 14243 20213
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 17218 20204 17224 20256
rect 17276 20204 17282 20256
rect 18598 20204 18604 20256
rect 18656 20244 18662 20256
rect 19061 20247 19119 20253
rect 19061 20244 19073 20247
rect 18656 20216 19073 20244
rect 18656 20204 18662 20216
rect 19061 20213 19073 20216
rect 19107 20213 19119 20247
rect 19061 20207 19119 20213
rect 20806 20204 20812 20256
rect 20864 20244 20870 20256
rect 20993 20247 21051 20253
rect 20993 20244 21005 20247
rect 20864 20216 21005 20244
rect 20864 20204 20870 20216
rect 20993 20213 21005 20216
rect 21039 20213 21051 20247
rect 20993 20207 21051 20213
rect 21174 20204 21180 20256
rect 21232 20204 21238 20256
rect 21450 20204 21456 20256
rect 21508 20244 21514 20256
rect 22066 20244 22094 20284
rect 22465 20281 22477 20284
rect 22511 20281 22523 20315
rect 22465 20275 22523 20281
rect 21508 20216 22094 20244
rect 21508 20204 21514 20216
rect 22278 20204 22284 20256
rect 22336 20204 22342 20256
rect 552 20154 23368 20176
rect 552 20102 19022 20154
rect 19074 20102 19086 20154
rect 19138 20102 19150 20154
rect 19202 20102 19214 20154
rect 19266 20102 19278 20154
rect 19330 20102 23368 20154
rect 552 20080 23368 20102
rect 5258 20040 5264 20052
rect 4448 20012 5264 20040
rect 4448 19913 4476 20012
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 5350 20000 5356 20052
rect 5408 20000 5414 20052
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 10100 20012 13032 20040
rect 10100 20000 10106 20012
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 4617 19907 4675 19913
rect 4617 19873 4629 19907
rect 4663 19904 4675 19907
rect 5261 19907 5319 19913
rect 5261 19904 5273 19907
rect 4663 19876 5273 19904
rect 4663 19873 4675 19876
rect 4617 19867 4675 19873
rect 5261 19873 5273 19876
rect 5307 19904 5319 19907
rect 5368 19904 5396 20000
rect 5629 19975 5687 19981
rect 5629 19941 5641 19975
rect 5675 19972 5687 19975
rect 9401 19975 9459 19981
rect 5675 19944 8800 19972
rect 5675 19941 5687 19944
rect 5629 19935 5687 19941
rect 6840 19916 6868 19944
rect 8772 19916 8800 19944
rect 9401 19941 9413 19975
rect 9447 19972 9459 19975
rect 10226 19972 10232 19984
rect 9447 19944 10232 19972
rect 9447 19941 9459 19944
rect 9401 19935 9459 19941
rect 10226 19932 10232 19944
rect 10284 19932 10290 19984
rect 11057 19975 11115 19981
rect 11057 19941 11069 19975
rect 11103 19972 11115 19975
rect 11330 19972 11336 19984
rect 11103 19944 11336 19972
rect 11103 19941 11115 19944
rect 11057 19935 11115 19941
rect 11330 19932 11336 19944
rect 11388 19932 11394 19984
rect 13004 19972 13032 20012
rect 13078 20000 13084 20052
rect 13136 20040 13142 20052
rect 13538 20040 13544 20052
rect 13136 20012 13544 20040
rect 13136 20000 13142 20012
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 17218 20000 17224 20052
rect 17276 20000 17282 20052
rect 17494 20000 17500 20052
rect 17552 20000 17558 20052
rect 18046 20040 18052 20052
rect 17604 20012 18052 20040
rect 13004 19944 13584 19972
rect 5307 19876 5396 19904
rect 5537 19907 5595 19913
rect 5307 19873 5319 19876
rect 5261 19867 5319 19873
rect 5537 19873 5549 19907
rect 5583 19904 5595 19907
rect 5718 19904 5724 19916
rect 5583 19876 5724 19904
rect 5583 19873 5595 19876
rect 5537 19867 5595 19873
rect 5718 19864 5724 19876
rect 5776 19904 5782 19916
rect 5905 19907 5963 19913
rect 5905 19904 5917 19907
rect 5776 19876 5917 19904
rect 5776 19864 5782 19876
rect 5905 19873 5917 19876
rect 5951 19873 5963 19907
rect 5905 19867 5963 19873
rect 6822 19864 6828 19916
rect 6880 19864 6886 19916
rect 7742 19864 7748 19916
rect 7800 19904 7806 19916
rect 8389 19907 8447 19913
rect 8389 19904 8401 19907
rect 7800 19876 8401 19904
rect 7800 19864 7806 19876
rect 8389 19873 8401 19876
rect 8435 19873 8447 19907
rect 8389 19867 8447 19873
rect 8754 19864 8760 19916
rect 8812 19864 8818 19916
rect 10042 19864 10048 19916
rect 10100 19864 10106 19916
rect 10244 19904 10272 19932
rect 10965 19907 11023 19913
rect 10965 19904 10977 19907
rect 10244 19876 10977 19904
rect 10965 19873 10977 19876
rect 11011 19873 11023 19907
rect 10965 19867 11023 19873
rect 11146 19864 11152 19916
rect 11204 19864 11210 19916
rect 11425 19907 11483 19913
rect 11425 19873 11437 19907
rect 11471 19873 11483 19907
rect 11425 19867 11483 19873
rect 4246 19796 4252 19848
rect 4304 19836 4310 19848
rect 4341 19839 4399 19845
rect 4341 19836 4353 19839
rect 4304 19808 4353 19836
rect 4304 19796 4310 19808
rect 4341 19805 4353 19808
rect 4387 19805 4399 19839
rect 4341 19799 4399 19805
rect 4890 19796 4896 19848
rect 4948 19836 4954 19848
rect 5166 19845 5172 19848
rect 5123 19839 5172 19845
rect 5123 19836 5135 19839
rect 4948 19808 5135 19836
rect 4948 19796 4954 19808
rect 5123 19805 5135 19808
rect 5169 19805 5172 19839
rect 5123 19799 5172 19805
rect 5166 19796 5172 19799
rect 5224 19796 5230 19848
rect 9766 19796 9772 19848
rect 9824 19796 9830 19848
rect 10689 19839 10747 19845
rect 10689 19805 10701 19839
rect 10735 19836 10747 19839
rect 11440 19836 11468 19867
rect 11606 19864 11612 19916
rect 11664 19864 11670 19916
rect 12713 19907 12771 19913
rect 12713 19904 12725 19907
rect 12098 19890 12725 19904
rect 12084 19876 12725 19890
rect 10735 19808 11468 19836
rect 11624 19836 11652 19864
rect 12084 19836 12112 19876
rect 12713 19873 12725 19876
rect 12759 19873 12771 19907
rect 12713 19867 12771 19873
rect 12805 19907 12863 19913
rect 12805 19873 12817 19907
rect 12851 19873 12863 19907
rect 12805 19867 12863 19873
rect 11624 19808 12112 19836
rect 10735 19805 10747 19808
rect 10689 19799 10747 19805
rect 4801 19771 4859 19777
rect 4801 19737 4813 19771
rect 4847 19768 4859 19771
rect 5258 19768 5264 19780
rect 4847 19740 5264 19768
rect 4847 19737 4859 19740
rect 4801 19731 4859 19737
rect 5258 19728 5264 19740
rect 5316 19728 5322 19780
rect 7098 19728 7104 19780
rect 7156 19728 7162 19780
rect 11440 19768 11468 19808
rect 12342 19796 12348 19848
rect 12400 19796 12406 19848
rect 12820 19768 12848 19867
rect 13354 19864 13360 19916
rect 13412 19904 13418 19916
rect 13449 19907 13507 19913
rect 13449 19904 13461 19907
rect 13412 19876 13461 19904
rect 13412 19864 13418 19876
rect 13449 19873 13461 19876
rect 13495 19873 13507 19907
rect 13449 19867 13507 19873
rect 13556 19845 13584 19944
rect 15948 19944 16896 19972
rect 13725 19907 13783 19913
rect 13725 19873 13737 19907
rect 13771 19904 13783 19907
rect 13817 19907 13875 19913
rect 13817 19904 13829 19907
rect 13771 19876 13829 19904
rect 13771 19873 13783 19876
rect 13725 19867 13783 19873
rect 13817 19873 13829 19876
rect 13863 19873 13875 19907
rect 14642 19904 14648 19916
rect 13817 19867 13875 19873
rect 13924 19876 14648 19904
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19836 13599 19839
rect 13924 19836 13952 19876
rect 14642 19864 14648 19876
rect 14700 19864 14706 19916
rect 15746 19864 15752 19916
rect 15804 19864 15810 19916
rect 15948 19913 15976 19944
rect 16868 19913 16896 19944
rect 15933 19907 15991 19913
rect 15933 19873 15945 19907
rect 15979 19873 15991 19907
rect 15933 19867 15991 19873
rect 16393 19907 16451 19913
rect 16393 19873 16405 19907
rect 16439 19873 16451 19907
rect 16393 19867 16451 19873
rect 16853 19907 16911 19913
rect 16853 19873 16865 19907
rect 16899 19904 16911 19907
rect 17236 19904 17264 20000
rect 17512 19913 17540 20000
rect 17604 19913 17632 20012
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 18230 20000 18236 20052
rect 18288 20000 18294 20052
rect 18598 20000 18604 20052
rect 18656 20000 18662 20052
rect 22002 20000 22008 20052
rect 22060 20000 22066 20052
rect 18248 19972 18276 20000
rect 17788 19944 18276 19972
rect 16899 19876 17264 19904
rect 17497 19907 17555 19913
rect 16899 19873 16911 19876
rect 16853 19867 16911 19873
rect 17497 19873 17509 19907
rect 17543 19873 17555 19907
rect 17497 19867 17555 19873
rect 17589 19907 17647 19913
rect 17589 19873 17601 19907
rect 17635 19873 17647 19907
rect 17589 19867 17647 19873
rect 13587 19808 13952 19836
rect 14001 19839 14059 19845
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 14001 19805 14013 19839
rect 14047 19805 14059 19839
rect 14001 19799 14059 19805
rect 14016 19768 14044 19799
rect 15194 19796 15200 19848
rect 15252 19836 15258 19848
rect 16408 19836 16436 19867
rect 15252 19808 16436 19836
rect 15252 19796 15258 19808
rect 17218 19796 17224 19848
rect 17276 19796 17282 19848
rect 11440 19740 12848 19768
rect 13832 19740 14044 19768
rect 15933 19771 15991 19777
rect 13832 19712 13860 19740
rect 15933 19737 15945 19771
rect 15979 19768 15991 19771
rect 17604 19768 17632 19867
rect 17788 19845 17816 19944
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19904 18291 19907
rect 18616 19904 18644 20000
rect 18690 19932 18696 19984
rect 18748 19972 18754 19984
rect 19061 19975 19119 19981
rect 19061 19972 19073 19975
rect 18748 19944 19073 19972
rect 18748 19932 18754 19944
rect 19061 19941 19073 19944
rect 19107 19941 19119 19975
rect 19061 19935 19119 19941
rect 19245 19975 19303 19981
rect 19245 19941 19257 19975
rect 19291 19972 19303 19975
rect 19291 19944 20024 19972
rect 19291 19941 19303 19944
rect 19245 19935 19303 19941
rect 18279 19876 18644 19904
rect 18877 19907 18935 19913
rect 18279 19873 18291 19876
rect 18233 19867 18291 19873
rect 18877 19873 18889 19907
rect 18923 19873 18935 19907
rect 18877 19867 18935 19873
rect 18969 19907 19027 19913
rect 18969 19873 18981 19907
rect 19015 19904 19027 19907
rect 19260 19904 19288 19935
rect 19996 19916 20024 19944
rect 19015 19876 19288 19904
rect 19337 19907 19395 19913
rect 19015 19873 19027 19876
rect 18969 19867 19027 19873
rect 19337 19873 19349 19907
rect 19383 19873 19395 19907
rect 19337 19867 19395 19873
rect 17773 19839 17831 19845
rect 17773 19805 17785 19839
rect 17819 19805 17831 19839
rect 17773 19799 17831 19805
rect 18049 19839 18107 19845
rect 18049 19805 18061 19839
rect 18095 19836 18107 19839
rect 18892 19836 18920 19867
rect 19352 19836 19380 19867
rect 19978 19864 19984 19916
rect 20036 19864 20042 19916
rect 20714 19864 20720 19916
rect 20772 19904 20778 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20772 19876 20913 19904
rect 20772 19864 20778 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 21266 19904 21272 19916
rect 21131 19876 21272 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 21266 19864 21272 19876
rect 21324 19904 21330 19916
rect 21542 19904 21548 19916
rect 21324 19876 21548 19904
rect 21324 19864 21330 19876
rect 21542 19864 21548 19876
rect 21600 19864 21606 19916
rect 21913 19907 21971 19913
rect 21913 19873 21925 19907
rect 21959 19904 21971 19907
rect 22020 19904 22048 20000
rect 21959 19876 22048 19904
rect 21959 19873 21971 19876
rect 21913 19867 21971 19873
rect 18095 19808 19380 19836
rect 18095 19805 18107 19808
rect 18049 19799 18107 19805
rect 15979 19740 17632 19768
rect 17681 19771 17739 19777
rect 15979 19737 15991 19740
rect 15933 19731 15991 19737
rect 17681 19737 17693 19771
rect 17727 19768 17739 19771
rect 18064 19768 18092 19799
rect 17727 19740 18092 19768
rect 17727 19737 17739 19740
rect 17681 19731 17739 19737
rect 4985 19703 5043 19709
rect 4985 19669 4997 19703
rect 5031 19700 5043 19703
rect 6914 19700 6920 19712
rect 5031 19672 6920 19700
rect 5031 19669 5043 19672
rect 4985 19663 5043 19669
rect 6914 19660 6920 19672
rect 6972 19660 6978 19712
rect 12526 19660 12532 19712
rect 12584 19660 12590 19712
rect 13814 19660 13820 19712
rect 13872 19660 13878 19712
rect 18414 19660 18420 19712
rect 18472 19660 18478 19712
rect 18690 19660 18696 19712
rect 18748 19660 18754 19712
rect 19150 19660 19156 19712
rect 19208 19660 19214 19712
rect 21082 19660 21088 19712
rect 21140 19660 21146 19712
rect 21821 19703 21879 19709
rect 21821 19669 21833 19703
rect 21867 19700 21879 19703
rect 22186 19700 22192 19712
rect 21867 19672 22192 19700
rect 21867 19669 21879 19672
rect 21821 19663 21879 19669
rect 22186 19660 22192 19672
rect 22244 19660 22250 19712
rect 552 19610 23368 19632
rect 552 19558 3662 19610
rect 3714 19558 3726 19610
rect 3778 19558 3790 19610
rect 3842 19558 3854 19610
rect 3906 19558 3918 19610
rect 3970 19558 23368 19610
rect 552 19536 23368 19558
rect 5350 19456 5356 19508
rect 5408 19456 5414 19508
rect 11425 19499 11483 19505
rect 11425 19465 11437 19499
rect 11471 19496 11483 19499
rect 12250 19496 12256 19508
rect 11471 19468 12256 19496
rect 11471 19465 11483 19468
rect 11425 19459 11483 19465
rect 5368 19360 5396 19456
rect 8205 19431 8263 19437
rect 8205 19397 8217 19431
rect 8251 19428 8263 19431
rect 9122 19428 9128 19440
rect 8251 19400 9128 19428
rect 8251 19397 8263 19400
rect 8205 19391 8263 19397
rect 9122 19388 9128 19400
rect 9180 19388 9186 19440
rect 5092 19332 5396 19360
rect 4430 19252 4436 19304
rect 4488 19252 4494 19304
rect 4801 19295 4859 19301
rect 4801 19261 4813 19295
rect 4847 19292 4859 19295
rect 4890 19292 4896 19304
rect 4847 19264 4896 19292
rect 4847 19261 4859 19264
rect 4801 19255 4859 19261
rect 4890 19252 4896 19264
rect 4948 19252 4954 19304
rect 5092 19301 5120 19332
rect 8386 19320 8392 19372
rect 8444 19360 8450 19372
rect 8444 19332 8892 19360
rect 8444 19320 8450 19332
rect 4985 19295 5043 19301
rect 4985 19261 4997 19295
rect 5031 19261 5043 19295
rect 4985 19255 5043 19261
rect 5077 19295 5135 19301
rect 5077 19261 5089 19295
rect 5123 19261 5135 19295
rect 5077 19255 5135 19261
rect 5353 19295 5411 19301
rect 5353 19261 5365 19295
rect 5399 19261 5411 19295
rect 5353 19255 5411 19261
rect 5629 19295 5687 19301
rect 5629 19261 5641 19295
rect 5675 19292 5687 19295
rect 5718 19292 5724 19304
rect 5675 19264 5724 19292
rect 5675 19261 5687 19264
rect 5629 19255 5687 19261
rect 4448 19224 4476 19252
rect 5000 19224 5028 19255
rect 4448 19196 5028 19224
rect 5368 19224 5396 19255
rect 5718 19252 5724 19264
rect 5776 19252 5782 19304
rect 5810 19252 5816 19304
rect 5868 19252 5874 19304
rect 5994 19252 6000 19304
rect 6052 19292 6058 19304
rect 6181 19295 6239 19301
rect 6181 19292 6193 19295
rect 6052 19264 6193 19292
rect 6052 19252 6058 19264
rect 6181 19261 6193 19264
rect 6227 19261 6239 19295
rect 6181 19255 6239 19261
rect 7098 19252 7104 19304
rect 7156 19252 7162 19304
rect 7282 19252 7288 19304
rect 7340 19292 7346 19304
rect 7377 19295 7435 19301
rect 7377 19292 7389 19295
rect 7340 19264 7389 19292
rect 7340 19252 7346 19264
rect 7377 19261 7389 19264
rect 7423 19261 7435 19295
rect 7377 19255 7435 19261
rect 8202 19252 8208 19304
rect 8260 19292 8266 19304
rect 8864 19301 8892 19332
rect 9766 19320 9772 19372
rect 9824 19320 9830 19372
rect 11146 19360 11152 19372
rect 10980 19332 11152 19360
rect 8757 19295 8815 19301
rect 8757 19292 8769 19295
rect 8260 19264 8769 19292
rect 8260 19252 8266 19264
rect 8757 19261 8769 19264
rect 8803 19261 8815 19295
rect 8757 19255 8815 19261
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19261 8907 19295
rect 8849 19255 8907 19261
rect 9033 19295 9091 19301
rect 9033 19261 9045 19295
rect 9079 19292 9091 19295
rect 9784 19292 9812 19320
rect 9079 19264 9812 19292
rect 9079 19261 9091 19264
rect 9033 19255 9091 19261
rect 10226 19252 10232 19304
rect 10284 19252 10290 19304
rect 10413 19295 10471 19301
rect 10413 19261 10425 19295
rect 10459 19292 10471 19295
rect 10980 19292 11008 19332
rect 11146 19320 11152 19332
rect 11204 19320 11210 19372
rect 11241 19363 11299 19369
rect 11241 19329 11253 19363
rect 11287 19360 11299 19363
rect 11440 19360 11468 19459
rect 12250 19456 12256 19468
rect 12308 19456 12314 19508
rect 15746 19456 15752 19508
rect 15804 19456 15810 19508
rect 18800 19468 19932 19496
rect 12526 19388 12532 19440
rect 12584 19428 12590 19440
rect 15473 19431 15531 19437
rect 15473 19428 15485 19431
rect 12584 19400 12664 19428
rect 12584 19388 12590 19400
rect 11287 19332 11468 19360
rect 11287 19329 11299 19332
rect 11241 19323 11299 19329
rect 11514 19320 11520 19372
rect 11572 19320 11578 19372
rect 11790 19320 11796 19372
rect 11848 19320 11854 19372
rect 12158 19320 12164 19372
rect 12216 19360 12222 19372
rect 12216 19332 12480 19360
rect 12636 19334 12664 19400
rect 14660 19400 15485 19428
rect 12216 19320 12222 19332
rect 10459 19264 11008 19292
rect 11333 19295 11391 19301
rect 10459 19261 10471 19264
rect 10413 19255 10471 19261
rect 11333 19261 11345 19295
rect 11379 19292 11391 19295
rect 11532 19292 11560 19320
rect 11379 19264 11560 19292
rect 11609 19295 11667 19301
rect 11379 19261 11391 19264
rect 11333 19255 11391 19261
rect 11609 19261 11621 19295
rect 11655 19261 11667 19295
rect 11609 19255 11667 19261
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19261 12311 19295
rect 12253 19255 12311 19261
rect 12345 19295 12403 19301
rect 12345 19261 12357 19295
rect 12391 19292 12403 19295
rect 12452 19292 12480 19332
rect 12544 19306 12664 19334
rect 13446 19320 13452 19372
rect 13504 19360 13510 19372
rect 13909 19363 13967 19369
rect 13504 19332 13768 19360
rect 13504 19320 13510 19332
rect 12544 19301 12572 19306
rect 12391 19264 12480 19292
rect 12509 19295 12572 19301
rect 12391 19261 12403 19264
rect 12345 19255 12403 19261
rect 12509 19261 12521 19295
rect 12555 19264 12572 19295
rect 13740 19292 13768 19332
rect 13909 19329 13921 19363
rect 13955 19329 13967 19363
rect 13909 19323 13967 19329
rect 13817 19295 13875 19301
rect 13817 19292 13829 19295
rect 13740 19264 13829 19292
rect 12555 19261 12567 19264
rect 12509 19255 12567 19261
rect 13817 19261 13829 19264
rect 13863 19261 13875 19295
rect 13817 19255 13875 19261
rect 6012 19224 6040 19252
rect 5368 19196 6040 19224
rect 6089 19227 6147 19233
rect 6089 19193 6101 19227
rect 6135 19224 6147 19227
rect 7300 19224 7328 19252
rect 10428 19224 10456 19255
rect 6135 19196 7328 19224
rect 8312 19196 10456 19224
rect 6135 19193 6147 19196
rect 6089 19187 6147 19193
rect 4706 19116 4712 19168
rect 4764 19156 4770 19168
rect 4801 19159 4859 19165
rect 4801 19156 4813 19159
rect 4764 19128 4813 19156
rect 4764 19116 4770 19128
rect 4801 19125 4813 19128
rect 4847 19125 4859 19159
rect 4801 19119 4859 19125
rect 4890 19116 4896 19168
rect 4948 19156 4954 19168
rect 5169 19159 5227 19165
rect 5169 19156 5181 19159
rect 4948 19128 5181 19156
rect 4948 19116 4954 19128
rect 5169 19125 5181 19128
rect 5215 19156 5227 19159
rect 5350 19156 5356 19168
rect 5215 19128 5356 19156
rect 5215 19125 5227 19128
rect 5169 19119 5227 19125
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 5534 19116 5540 19168
rect 5592 19116 5598 19168
rect 6914 19116 6920 19168
rect 6972 19156 6978 19168
rect 8312 19156 8340 19196
rect 10502 19184 10508 19236
rect 10560 19224 10566 19236
rect 11348 19224 11376 19255
rect 10560 19196 11376 19224
rect 10560 19184 10566 19196
rect 11422 19184 11428 19236
rect 11480 19224 11486 19236
rect 11624 19224 11652 19255
rect 11480 19196 11652 19224
rect 12268 19224 12296 19255
rect 13924 19224 13952 19323
rect 13998 19320 14004 19372
rect 14056 19320 14062 19372
rect 14090 19320 14096 19372
rect 14148 19360 14154 19372
rect 14553 19363 14611 19369
rect 14553 19360 14565 19363
rect 14148 19332 14565 19360
rect 14148 19320 14154 19332
rect 14553 19329 14565 19332
rect 14599 19329 14611 19363
rect 14553 19323 14611 19329
rect 14016 19292 14044 19320
rect 14660 19292 14688 19400
rect 15473 19397 15485 19400
rect 15519 19428 15531 19431
rect 15764 19428 15792 19456
rect 15519 19400 15792 19428
rect 15519 19397 15531 19400
rect 15473 19391 15531 19397
rect 17218 19388 17224 19440
rect 17276 19428 17282 19440
rect 18141 19431 18199 19437
rect 18141 19428 18153 19431
rect 17276 19400 18153 19428
rect 17276 19388 17282 19400
rect 16666 19320 16672 19372
rect 16724 19320 16730 19372
rect 14016 19264 14688 19292
rect 15378 19252 15384 19304
rect 15436 19252 15442 19304
rect 16298 19252 16304 19304
rect 16356 19252 16362 19304
rect 16684 19292 16712 19320
rect 17604 19301 17632 19400
rect 18141 19397 18153 19400
rect 18187 19397 18199 19431
rect 18141 19391 18199 19397
rect 18414 19320 18420 19372
rect 18472 19360 18478 19372
rect 18800 19360 18828 19468
rect 18874 19388 18880 19440
rect 18932 19428 18938 19440
rect 19150 19428 19156 19440
rect 18932 19400 19156 19428
rect 18932 19388 18938 19400
rect 19150 19388 19156 19400
rect 19208 19428 19214 19440
rect 19429 19431 19487 19437
rect 19429 19428 19441 19431
rect 19208 19400 19441 19428
rect 19208 19388 19214 19400
rect 19429 19397 19441 19400
rect 19475 19397 19487 19431
rect 19429 19391 19487 19397
rect 18969 19363 19027 19369
rect 18969 19360 18981 19363
rect 18472 19332 18981 19360
rect 18472 19320 18478 19332
rect 18969 19329 18981 19332
rect 19015 19329 19027 19363
rect 19904 19360 19932 19468
rect 19978 19456 19984 19508
rect 20036 19456 20042 19508
rect 21174 19456 21180 19508
rect 21232 19496 21238 19508
rect 21361 19499 21419 19505
rect 21361 19496 21373 19499
rect 21232 19468 21373 19496
rect 21232 19456 21238 19468
rect 21361 19465 21373 19468
rect 21407 19465 21419 19499
rect 21361 19459 21419 19465
rect 21450 19456 21456 19508
rect 21508 19456 21514 19508
rect 21634 19456 21640 19508
rect 21692 19496 21698 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21692 19468 22017 19496
rect 21692 19456 21698 19468
rect 22005 19465 22017 19468
rect 22051 19496 22063 19499
rect 22051 19468 22416 19496
rect 22051 19465 22063 19468
rect 22005 19459 22063 19465
rect 21468 19428 21496 19456
rect 20640 19400 21496 19428
rect 20533 19363 20591 19369
rect 18969 19323 19027 19329
rect 19168 19332 19840 19360
rect 19904 19332 20024 19360
rect 17221 19295 17279 19301
rect 17221 19292 17233 19295
rect 16684 19264 17233 19292
rect 17221 19261 17233 19264
rect 17267 19261 17279 19295
rect 17221 19255 17279 19261
rect 17589 19295 17647 19301
rect 17589 19261 17601 19295
rect 17635 19261 17647 19295
rect 17589 19255 17647 19261
rect 12268 19196 13952 19224
rect 17236 19224 17264 19255
rect 17678 19252 17684 19304
rect 17736 19292 17742 19304
rect 19061 19295 19119 19301
rect 19061 19292 19073 19295
rect 17736 19264 19073 19292
rect 17736 19252 17742 19264
rect 19061 19261 19073 19264
rect 19107 19292 19119 19295
rect 19168 19292 19196 19332
rect 19107 19264 19196 19292
rect 19812 19292 19840 19332
rect 19889 19295 19947 19301
rect 19889 19292 19901 19295
rect 19812 19264 19901 19292
rect 19107 19261 19119 19264
rect 19061 19255 19119 19261
rect 19889 19261 19901 19264
rect 19935 19261 19947 19295
rect 19996 19292 20024 19332
rect 20533 19329 20545 19363
rect 20579 19360 20591 19363
rect 20640 19360 20668 19400
rect 20579 19332 20668 19360
rect 20579 19329 20591 19332
rect 20533 19323 20591 19329
rect 20640 19304 20668 19332
rect 20732 19332 21036 19360
rect 20732 19304 20760 19332
rect 20073 19295 20131 19301
rect 20073 19292 20085 19295
rect 19996 19264 20085 19292
rect 19889 19255 19947 19261
rect 20073 19261 20085 19264
rect 20119 19261 20131 19295
rect 20073 19255 20131 19261
rect 20257 19295 20315 19301
rect 20257 19261 20269 19295
rect 20303 19261 20315 19295
rect 20257 19255 20315 19261
rect 18509 19227 18567 19233
rect 18509 19224 18521 19227
rect 17236 19196 18521 19224
rect 11480 19184 11486 19196
rect 12406 19168 12434 19196
rect 18509 19193 18521 19196
rect 18555 19193 18567 19227
rect 18509 19187 18567 19193
rect 18782 19184 18788 19236
rect 18840 19224 18846 19236
rect 19797 19227 19855 19233
rect 19797 19224 19809 19227
rect 18840 19196 19809 19224
rect 18840 19184 18846 19196
rect 19797 19193 19809 19196
rect 19843 19193 19855 19227
rect 19797 19187 19855 19193
rect 6972 19128 8340 19156
rect 6972 19116 6978 19128
rect 8386 19116 8392 19168
rect 8444 19116 8450 19168
rect 12342 19116 12348 19168
rect 12400 19128 12434 19168
rect 12400 19116 12406 19128
rect 12710 19116 12716 19168
rect 12768 19116 12774 19168
rect 16853 19159 16911 19165
rect 16853 19125 16865 19159
rect 16899 19156 16911 19159
rect 17310 19156 17316 19168
rect 16899 19128 17316 19156
rect 16899 19125 16911 19128
rect 16853 19119 16911 19125
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 18046 19116 18052 19168
rect 18104 19116 18110 19168
rect 18598 19116 18604 19168
rect 18656 19156 18662 19168
rect 18693 19159 18751 19165
rect 18693 19156 18705 19159
rect 18656 19128 18705 19156
rect 18656 19116 18662 19128
rect 18693 19125 18705 19128
rect 18739 19125 18751 19159
rect 18693 19119 18751 19125
rect 19337 19159 19395 19165
rect 19337 19125 19349 19159
rect 19383 19156 19395 19159
rect 19518 19156 19524 19168
rect 19383 19128 19524 19156
rect 19383 19125 19395 19128
rect 19337 19119 19395 19125
rect 19518 19116 19524 19128
rect 19576 19116 19582 19168
rect 20272 19156 20300 19255
rect 20346 19252 20352 19304
rect 20404 19252 20410 19304
rect 20622 19252 20628 19304
rect 20680 19252 20686 19304
rect 20714 19252 20720 19304
rect 20772 19252 20778 19304
rect 20806 19252 20812 19304
rect 20864 19252 20870 19304
rect 21008 19301 21036 19332
rect 21082 19320 21088 19372
rect 21140 19360 21146 19372
rect 21453 19363 21511 19369
rect 21453 19360 21465 19363
rect 21140 19332 21465 19360
rect 21140 19320 21146 19332
rect 21453 19329 21465 19332
rect 21499 19329 21511 19363
rect 21453 19323 21511 19329
rect 21358 19301 21364 19304
rect 20901 19295 20959 19301
rect 20901 19261 20913 19295
rect 20947 19261 20959 19295
rect 20901 19255 20959 19261
rect 20993 19295 21051 19301
rect 20993 19261 21005 19295
rect 21039 19261 21051 19295
rect 21349 19295 21364 19301
rect 21349 19292 21361 19295
rect 20993 19255 21051 19261
rect 21284 19264 21361 19292
rect 20364 19224 20392 19252
rect 20916 19224 20944 19255
rect 21284 19233 21312 19264
rect 21349 19261 21361 19264
rect 21349 19255 21364 19261
rect 21358 19252 21364 19255
rect 21416 19252 21422 19304
rect 22278 19292 22284 19304
rect 22112 19264 22284 19292
rect 20364 19196 20944 19224
rect 21269 19227 21327 19233
rect 21269 19193 21281 19227
rect 21315 19193 21327 19227
rect 21269 19187 21327 19193
rect 21989 19227 22047 19233
rect 21989 19193 22001 19227
rect 22035 19224 22047 19227
rect 22112 19224 22140 19264
rect 22278 19252 22284 19264
rect 22336 19252 22342 19304
rect 22388 19292 22416 19468
rect 22557 19295 22615 19301
rect 22557 19292 22569 19295
rect 22388 19264 22569 19292
rect 22557 19261 22569 19264
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 22035 19196 22140 19224
rect 22035 19193 22047 19196
rect 21989 19187 22047 19193
rect 22186 19184 22192 19236
rect 22244 19224 22250 19236
rect 22465 19227 22523 19233
rect 22465 19224 22477 19227
rect 22244 19196 22477 19224
rect 22244 19184 22250 19196
rect 22465 19193 22477 19196
rect 22511 19193 22523 19227
rect 22465 19187 22523 19193
rect 20438 19156 20444 19168
rect 20272 19128 20444 19156
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 20533 19159 20591 19165
rect 20533 19125 20545 19159
rect 20579 19156 20591 19159
rect 20714 19156 20720 19168
rect 20579 19128 20720 19156
rect 20579 19125 20591 19128
rect 20533 19119 20591 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 20990 19116 20996 19168
rect 21048 19156 21054 19168
rect 21729 19159 21787 19165
rect 21729 19156 21741 19159
rect 21048 19128 21741 19156
rect 21048 19116 21054 19128
rect 21729 19125 21741 19128
rect 21775 19125 21787 19159
rect 21729 19119 21787 19125
rect 21818 19116 21824 19168
rect 21876 19116 21882 19168
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22379 19159 22437 19165
rect 22379 19156 22391 19159
rect 22152 19128 22391 19156
rect 22152 19116 22158 19128
rect 22379 19125 22391 19128
rect 22425 19125 22437 19159
rect 22379 19119 22437 19125
rect 552 19066 23368 19088
rect 552 19014 19022 19066
rect 19074 19014 19086 19066
rect 19138 19014 19150 19066
rect 19202 19014 19214 19066
rect 19266 19014 19278 19066
rect 19330 19014 23368 19066
rect 552 18992 23368 19014
rect 5534 18912 5540 18964
rect 5592 18912 5598 18964
rect 5718 18912 5724 18964
rect 5776 18952 5782 18964
rect 7926 18952 7932 18964
rect 5776 18924 7932 18952
rect 5776 18912 5782 18924
rect 7926 18912 7932 18924
rect 7984 18912 7990 18964
rect 8021 18955 8079 18961
rect 8021 18921 8033 18955
rect 8067 18952 8079 18955
rect 8386 18952 8392 18964
rect 8067 18924 8392 18952
rect 8067 18921 8079 18924
rect 8021 18915 8079 18921
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 9309 18955 9367 18961
rect 9309 18952 9321 18955
rect 9048 18924 9321 18952
rect 5552 18884 5580 18912
rect 5552 18856 7880 18884
rect 4706 18776 4712 18828
rect 4764 18816 4770 18828
rect 6181 18819 6239 18825
rect 6181 18816 6193 18819
rect 4764 18788 6193 18816
rect 4764 18776 4770 18788
rect 6181 18785 6193 18788
rect 6227 18785 6239 18819
rect 6181 18779 6239 18785
rect 6270 18776 6276 18828
rect 6328 18776 6334 18828
rect 6656 18825 6684 18856
rect 6641 18819 6699 18825
rect 6641 18785 6653 18819
rect 6687 18785 6699 18819
rect 6641 18779 6699 18785
rect 6822 18776 6828 18828
rect 6880 18776 6886 18828
rect 7852 18825 7880 18856
rect 7837 18819 7895 18825
rect 7837 18785 7849 18819
rect 7883 18785 7895 18819
rect 7944 18816 7972 18912
rect 8294 18844 8300 18896
rect 8352 18844 8358 18896
rect 8404 18884 8432 18912
rect 8481 18887 8539 18893
rect 8481 18884 8493 18887
rect 8404 18856 8493 18884
rect 8481 18853 8493 18856
rect 8527 18853 8539 18887
rect 8481 18847 8539 18853
rect 8021 18819 8079 18825
rect 8021 18816 8033 18819
rect 7944 18788 8033 18816
rect 7837 18779 7895 18785
rect 8021 18785 8033 18788
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 8202 18776 8208 18828
rect 8260 18776 8266 18828
rect 8312 18816 8340 18844
rect 8389 18819 8447 18825
rect 8389 18816 8401 18819
rect 8312 18788 8401 18816
rect 8389 18785 8401 18788
rect 8435 18785 8447 18819
rect 8389 18779 8447 18785
rect 8573 18819 8631 18825
rect 8573 18785 8585 18819
rect 8619 18816 8631 18819
rect 8754 18816 8760 18828
rect 8619 18788 8760 18816
rect 8619 18785 8631 18788
rect 8573 18779 8631 18785
rect 8754 18776 8760 18788
rect 8812 18816 8818 18828
rect 9048 18816 9076 18924
rect 9309 18921 9321 18924
rect 9355 18952 9367 18955
rect 10042 18952 10048 18964
rect 9355 18924 10048 18952
rect 9355 18921 9367 18924
rect 9309 18915 9367 18921
rect 10042 18912 10048 18924
rect 10100 18912 10106 18964
rect 10870 18912 10876 18964
rect 10928 18952 10934 18964
rect 15194 18952 15200 18964
rect 10928 18924 15200 18952
rect 10928 18912 10934 18924
rect 9122 18844 9128 18896
rect 9180 18884 9186 18896
rect 9180 18856 9996 18884
rect 9180 18844 9186 18856
rect 9232 18825 9260 18856
rect 8812 18788 9076 18816
rect 9217 18819 9275 18825
rect 8812 18776 8818 18788
rect 9217 18785 9229 18819
rect 9263 18785 9275 18819
rect 9217 18779 9275 18785
rect 9398 18776 9404 18828
rect 9456 18816 9462 18828
rect 9968 18825 9996 18856
rect 10704 18856 12388 18884
rect 9493 18819 9551 18825
rect 9493 18816 9505 18819
rect 9456 18788 9505 18816
rect 9456 18776 9462 18788
rect 9493 18785 9505 18788
rect 9539 18785 9551 18819
rect 9493 18779 9551 18785
rect 9953 18819 10011 18825
rect 9953 18785 9965 18819
rect 9999 18785 10011 18819
rect 9953 18779 10011 18785
rect 10413 18819 10471 18825
rect 10413 18785 10425 18819
rect 10459 18816 10471 18819
rect 10502 18816 10508 18828
rect 10459 18788 10508 18816
rect 10459 18785 10471 18788
rect 10413 18779 10471 18785
rect 5813 18751 5871 18757
rect 5813 18717 5825 18751
rect 5859 18717 5871 18751
rect 5813 18711 5871 18717
rect 5905 18751 5963 18757
rect 5905 18717 5917 18751
rect 5951 18748 5963 18751
rect 5994 18748 6000 18760
rect 5951 18720 6000 18748
rect 5951 18717 5963 18720
rect 5905 18711 5963 18717
rect 5828 18680 5856 18711
rect 5994 18708 6000 18720
rect 6052 18708 6058 18760
rect 6840 18680 6868 18776
rect 7653 18751 7711 18757
rect 7653 18717 7665 18751
rect 7699 18748 7711 18751
rect 8220 18748 8248 18776
rect 7699 18720 8248 18748
rect 7699 18717 7711 18720
rect 7653 18711 7711 18717
rect 5828 18652 6868 18680
rect 7852 18624 7880 18720
rect 9858 18708 9864 18760
rect 9916 18748 9922 18760
rect 10428 18748 10456 18779
rect 10502 18776 10508 18788
rect 10560 18776 10566 18828
rect 9916 18720 10456 18748
rect 9916 18708 9922 18720
rect 8757 18683 8815 18689
rect 8757 18649 8769 18683
rect 8803 18680 8815 18683
rect 10704 18680 10732 18856
rect 12360 18825 12388 18856
rect 10781 18819 10839 18825
rect 10781 18785 10793 18819
rect 10827 18816 10839 18819
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 10827 18788 11437 18816
rect 10827 18785 10839 18788
rect 10781 18779 10839 18785
rect 11425 18785 11437 18788
rect 11471 18816 11483 18819
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 11471 18788 12173 18816
rect 11471 18785 11483 18788
rect 11425 18779 11483 18785
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12161 18779 12219 18785
rect 12345 18819 12403 18825
rect 12345 18785 12357 18819
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 13449 18819 13507 18825
rect 13449 18785 13461 18819
rect 13495 18785 13507 18819
rect 13556 18816 13584 18924
rect 15194 18912 15200 18924
rect 15252 18912 15258 18964
rect 18046 18912 18052 18964
rect 18104 18912 18110 18964
rect 18598 18912 18604 18964
rect 18656 18952 18662 18964
rect 19150 18952 19156 18964
rect 18656 18924 19156 18952
rect 18656 18912 18662 18924
rect 17589 18887 17647 18893
rect 17589 18884 17601 18887
rect 16500 18856 17601 18884
rect 16500 18828 16528 18856
rect 17589 18853 17601 18856
rect 17635 18884 17647 18887
rect 17678 18884 17684 18896
rect 17635 18856 17684 18884
rect 17635 18853 17647 18856
rect 17589 18847 17647 18853
rect 17678 18844 17684 18856
rect 17736 18844 17742 18896
rect 17773 18887 17831 18893
rect 17773 18853 17785 18887
rect 17819 18884 17831 18887
rect 18064 18884 18092 18912
rect 17819 18856 18092 18884
rect 17819 18853 17831 18856
rect 17773 18847 17831 18853
rect 13633 18819 13691 18825
rect 13633 18816 13645 18819
rect 13556 18788 13645 18816
rect 13449 18779 13507 18785
rect 13633 18785 13645 18788
rect 13679 18785 13691 18819
rect 13633 18779 13691 18785
rect 14461 18819 14519 18825
rect 14461 18785 14473 18819
rect 14507 18816 14519 18819
rect 14734 18816 14740 18828
rect 14507 18788 14740 18816
rect 14507 18785 14519 18788
rect 14461 18779 14519 18785
rect 11149 18751 11207 18757
rect 11149 18717 11161 18751
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18717 12127 18751
rect 12069 18711 12127 18717
rect 11164 18680 11192 18711
rect 8803 18652 11192 18680
rect 8803 18649 8815 18652
rect 8757 18643 8815 18649
rect 11790 18640 11796 18692
rect 11848 18680 11854 18692
rect 12084 18680 12112 18711
rect 12250 18708 12256 18760
rect 12308 18748 12314 18760
rect 13464 18748 13492 18779
rect 14734 18776 14740 18788
rect 14792 18816 14798 18828
rect 14829 18819 14887 18825
rect 14829 18816 14841 18819
rect 14792 18788 14841 18816
rect 14792 18776 14798 18788
rect 14829 18785 14841 18788
rect 14875 18785 14887 18819
rect 14829 18779 14887 18785
rect 14918 18776 14924 18828
rect 14976 18816 14982 18828
rect 15105 18819 15163 18825
rect 15105 18816 15117 18819
rect 14976 18788 15117 18816
rect 14976 18776 14982 18788
rect 15105 18785 15117 18788
rect 15151 18785 15163 18819
rect 15105 18779 15163 18785
rect 16482 18776 16488 18828
rect 16540 18776 16546 18828
rect 17497 18819 17555 18825
rect 17497 18816 17509 18819
rect 17328 18788 17509 18816
rect 17328 18760 17356 18788
rect 17497 18785 17509 18788
rect 17543 18785 17555 18819
rect 17497 18779 17555 18785
rect 18509 18819 18567 18825
rect 18509 18785 18521 18819
rect 18555 18816 18567 18819
rect 18708 18816 18736 18924
rect 19150 18912 19156 18924
rect 19208 18912 19214 18964
rect 19288 18912 19294 18964
rect 19346 18912 19352 18964
rect 19429 18955 19487 18961
rect 19429 18921 19441 18955
rect 19475 18952 19487 18955
rect 20346 18952 20352 18964
rect 19475 18924 20352 18952
rect 19475 18921 19487 18924
rect 19429 18915 19487 18921
rect 20346 18912 20352 18924
rect 20404 18912 20410 18964
rect 21174 18912 21180 18964
rect 21232 18912 21238 18964
rect 22465 18955 22523 18961
rect 22465 18921 22477 18955
rect 22511 18952 22523 18955
rect 22554 18952 22560 18964
rect 22511 18924 22560 18952
rect 22511 18921 22523 18924
rect 22465 18915 22523 18921
rect 22554 18912 22560 18924
rect 22612 18912 22618 18964
rect 19306 18884 19334 18912
rect 19306 18856 19748 18884
rect 18555 18788 18736 18816
rect 18555 18785 18567 18788
rect 18509 18779 18567 18785
rect 18782 18776 18788 18828
rect 18840 18816 18846 18828
rect 19061 18822 19119 18825
rect 18892 18819 19119 18822
rect 18892 18816 19073 18819
rect 18840 18794 19073 18816
rect 18840 18788 18920 18794
rect 18840 18776 18846 18788
rect 19061 18785 19073 18794
rect 19107 18785 19119 18819
rect 19061 18779 19119 18785
rect 19150 18776 19156 18828
rect 19208 18825 19214 18828
rect 19208 18819 19243 18825
rect 19231 18785 19243 18819
rect 19208 18779 19243 18785
rect 19208 18776 19214 18779
rect 19288 18776 19294 18828
rect 19346 18816 19352 18828
rect 19720 18825 19748 18856
rect 19521 18819 19579 18825
rect 19521 18816 19533 18819
rect 19346 18788 19533 18816
rect 19346 18776 19352 18788
rect 19521 18785 19533 18788
rect 19567 18785 19579 18819
rect 19521 18779 19579 18785
rect 19705 18819 19763 18825
rect 19705 18785 19717 18819
rect 19751 18785 19763 18819
rect 20364 18816 20392 18912
rect 20809 18819 20867 18825
rect 20809 18816 20821 18819
rect 20364 18788 20821 18816
rect 19705 18779 19763 18785
rect 20809 18785 20821 18788
rect 20855 18785 20867 18819
rect 21192 18816 21220 18912
rect 21269 18819 21327 18825
rect 21269 18816 21281 18819
rect 21192 18788 21281 18816
rect 20809 18779 20867 18785
rect 21269 18785 21281 18788
rect 21315 18785 21327 18819
rect 21269 18779 21327 18785
rect 21358 18776 21364 18828
rect 21416 18776 21422 18828
rect 22186 18776 22192 18828
rect 22244 18776 22250 18828
rect 12308 18720 13492 18748
rect 15657 18751 15715 18757
rect 12308 18708 12314 18720
rect 15657 18717 15669 18751
rect 15703 18748 15715 18751
rect 16390 18748 16396 18760
rect 15703 18720 16396 18748
rect 15703 18717 15715 18720
rect 15657 18711 15715 18717
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 17310 18708 17316 18760
rect 17368 18708 17374 18760
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18717 18659 18751
rect 18957 18751 19015 18757
rect 18957 18748 18969 18751
rect 18601 18711 18659 18717
rect 18892 18720 18969 18748
rect 12434 18680 12440 18692
rect 11848 18652 12440 18680
rect 11848 18640 11854 18652
rect 12434 18640 12440 18652
rect 12492 18640 12498 18692
rect 17773 18683 17831 18689
rect 17773 18649 17785 18683
rect 17819 18649 17831 18683
rect 17773 18643 17831 18649
rect 18616 18680 18644 18711
rect 18690 18680 18696 18692
rect 18616 18652 18696 18680
rect 6454 18572 6460 18624
rect 6512 18572 6518 18624
rect 7834 18572 7840 18624
rect 7892 18572 7898 18624
rect 9490 18572 9496 18624
rect 9548 18572 9554 18624
rect 12250 18572 12256 18624
rect 12308 18572 12314 18624
rect 12342 18572 12348 18624
rect 12400 18612 12406 18624
rect 13078 18612 13084 18624
rect 12400 18584 13084 18612
rect 12400 18572 12406 18584
rect 13078 18572 13084 18584
rect 13136 18572 13142 18624
rect 17788 18612 17816 18643
rect 18616 18612 18644 18652
rect 18690 18640 18696 18652
rect 18748 18640 18754 18692
rect 17788 18584 18644 18612
rect 18782 18572 18788 18624
rect 18840 18572 18846 18624
rect 18892 18612 18920 18720
rect 18957 18717 18969 18720
rect 19003 18717 19015 18751
rect 19426 18748 19432 18760
rect 18957 18711 19015 18717
rect 19306 18720 19432 18748
rect 18966 18612 18972 18624
rect 18892 18584 18972 18612
rect 18966 18572 18972 18584
rect 19024 18572 19030 18624
rect 19150 18572 19156 18624
rect 19208 18612 19214 18624
rect 19306 18612 19334 18720
rect 19426 18708 19432 18720
rect 19484 18748 19490 18760
rect 19484 18720 19564 18748
rect 19484 18708 19490 18720
rect 19536 18689 19564 18720
rect 20622 18708 20628 18760
rect 20680 18748 20686 18760
rect 20717 18751 20775 18757
rect 20717 18748 20729 18751
rect 20680 18720 20729 18748
rect 20680 18708 20686 18720
rect 20717 18717 20729 18720
rect 20763 18717 20775 18751
rect 20717 18711 20775 18717
rect 21082 18708 21088 18760
rect 21140 18748 21146 18760
rect 21545 18751 21603 18757
rect 21545 18748 21557 18751
rect 21140 18720 21557 18748
rect 21140 18708 21146 18720
rect 21545 18717 21557 18720
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 19521 18683 19579 18689
rect 19521 18649 19533 18683
rect 19567 18649 19579 18683
rect 19521 18643 19579 18649
rect 19208 18584 19334 18612
rect 19208 18572 19214 18584
rect 20438 18572 20444 18624
rect 20496 18572 20502 18624
rect 20622 18572 20628 18624
rect 20680 18572 20686 18624
rect 21358 18572 21364 18624
rect 21416 18612 21422 18624
rect 21453 18615 21511 18621
rect 21453 18612 21465 18615
rect 21416 18584 21465 18612
rect 21416 18572 21422 18584
rect 21453 18581 21465 18584
rect 21499 18581 21511 18615
rect 21453 18575 21511 18581
rect 552 18522 23368 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 23368 18522
rect 552 18448 23368 18470
rect 6086 18368 6092 18420
rect 6144 18368 6150 18420
rect 6365 18411 6423 18417
rect 6365 18377 6377 18411
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 6104 18340 6132 18368
rect 4172 18312 5396 18340
rect 4172 18281 4200 18312
rect 5368 18284 5396 18312
rect 5644 18312 6132 18340
rect 6380 18340 6408 18371
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 6972 18380 7788 18408
rect 6972 18368 6978 18380
rect 6380 18312 7052 18340
rect 4157 18275 4215 18281
rect 4157 18241 4169 18275
rect 4203 18241 4215 18275
rect 4157 18235 4215 18241
rect 4433 18275 4491 18281
rect 4433 18241 4445 18275
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18272 5043 18275
rect 5258 18272 5264 18284
rect 5031 18244 5264 18272
rect 5031 18241 5043 18244
rect 4985 18235 5043 18241
rect 4065 18207 4123 18213
rect 4065 18173 4077 18207
rect 4111 18204 4123 18207
rect 4246 18204 4252 18216
rect 4111 18176 4252 18204
rect 4111 18173 4123 18176
rect 4065 18167 4123 18173
rect 4246 18164 4252 18176
rect 4304 18164 4310 18216
rect 4448 18068 4476 18235
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 5350 18232 5356 18284
rect 5408 18232 5414 18284
rect 5644 18204 5672 18312
rect 5994 18232 6000 18284
rect 6052 18232 6058 18284
rect 6196 18244 6776 18272
rect 5474 18176 5672 18204
rect 5718 18164 5724 18216
rect 5776 18204 5782 18216
rect 6089 18207 6147 18213
rect 6089 18204 6101 18207
rect 5776 18176 6101 18204
rect 5776 18164 5782 18176
rect 6089 18173 6101 18176
rect 6135 18173 6147 18207
rect 6089 18167 6147 18173
rect 5810 18096 5816 18148
rect 5868 18136 5874 18148
rect 6196 18136 6224 18244
rect 6454 18164 6460 18216
rect 6512 18206 6518 18216
rect 6748 18213 6776 18244
rect 6914 18232 6920 18284
rect 6972 18232 6978 18284
rect 7024 18281 7052 18312
rect 7760 18281 7788 18380
rect 8754 18368 8760 18420
rect 8812 18368 8818 18420
rect 11790 18368 11796 18420
rect 11848 18368 11854 18420
rect 14734 18368 14740 18420
rect 14792 18368 14798 18420
rect 14829 18411 14887 18417
rect 14829 18377 14841 18411
rect 14875 18408 14887 18411
rect 14918 18408 14924 18420
rect 14875 18380 14924 18408
rect 14875 18377 14887 18380
rect 14829 18371 14887 18377
rect 7009 18275 7067 18281
rect 7009 18241 7021 18275
rect 7055 18272 7067 18275
rect 7745 18275 7803 18281
rect 7055 18244 7696 18272
rect 7055 18241 7067 18244
rect 7009 18235 7067 18241
rect 6549 18207 6607 18213
rect 6549 18206 6561 18207
rect 6512 18178 6561 18206
rect 6512 18164 6518 18178
rect 6549 18173 6561 18178
rect 6595 18173 6607 18207
rect 6549 18167 6607 18173
rect 6733 18207 6791 18213
rect 6733 18173 6745 18207
rect 6779 18173 6791 18207
rect 6932 18204 6960 18232
rect 7668 18213 7696 18244
rect 7745 18241 7757 18275
rect 7791 18241 7803 18275
rect 7745 18235 7803 18241
rect 8021 18275 8079 18281
rect 8021 18241 8033 18275
rect 8067 18272 8079 18275
rect 8202 18272 8208 18284
rect 8067 18244 8208 18272
rect 8067 18241 8079 18244
rect 8021 18235 8079 18241
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 8772 18213 8800 18368
rect 13078 18340 13084 18352
rect 12544 18312 13084 18340
rect 8849 18275 8907 18281
rect 8849 18241 8861 18275
rect 8895 18272 8907 18275
rect 9122 18272 9128 18284
rect 8895 18244 9128 18272
rect 8895 18241 8907 18244
rect 8849 18235 8907 18241
rect 9122 18232 9128 18244
rect 9180 18272 9186 18284
rect 9180 18244 10732 18272
rect 9180 18232 9186 18244
rect 7193 18207 7251 18213
rect 7193 18204 7205 18207
rect 6932 18176 7205 18204
rect 6733 18167 6791 18173
rect 7193 18173 7205 18176
rect 7239 18173 7251 18207
rect 7193 18167 7251 18173
rect 7653 18207 7711 18213
rect 7653 18173 7665 18207
rect 7699 18173 7711 18207
rect 7653 18167 7711 18173
rect 8757 18207 8815 18213
rect 8757 18173 8769 18207
rect 8803 18173 8815 18207
rect 8757 18167 8815 18173
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 10704 18213 10732 18244
rect 10870 18232 10876 18284
rect 10928 18232 10934 18284
rect 11701 18275 11759 18281
rect 11701 18241 11713 18275
rect 11747 18241 11759 18275
rect 12250 18272 12256 18284
rect 11701 18235 11759 18241
rect 11992 18244 12256 18272
rect 10321 18207 10379 18213
rect 10321 18204 10333 18207
rect 9456 18176 10333 18204
rect 9456 18164 9462 18176
rect 10321 18173 10333 18176
rect 10367 18173 10379 18207
rect 10321 18167 10379 18173
rect 10689 18207 10747 18213
rect 10689 18173 10701 18207
rect 10735 18173 10747 18207
rect 10689 18167 10747 18173
rect 5868 18108 6224 18136
rect 6641 18139 6699 18145
rect 5868 18096 5874 18108
rect 6641 18105 6653 18139
rect 6687 18136 6699 18139
rect 8294 18136 8300 18148
rect 6687 18108 8300 18136
rect 6687 18105 6699 18108
rect 6641 18099 6699 18105
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 10962 18096 10968 18148
rect 11020 18136 11026 18148
rect 11716 18136 11744 18235
rect 11992 18213 12020 18244
rect 12250 18232 12256 18244
rect 12308 18232 12314 18284
rect 12544 18281 12572 18312
rect 13078 18300 13084 18312
rect 13136 18300 13142 18352
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 12710 18232 12716 18284
rect 12768 18272 12774 18284
rect 12768 18244 13584 18272
rect 12768 18232 12774 18244
rect 12440 18216 12492 18222
rect 13556 18216 13584 18244
rect 11977 18207 12035 18213
rect 11977 18173 11989 18207
rect 12023 18173 12035 18207
rect 11977 18167 12035 18173
rect 12158 18164 12164 18216
rect 12216 18164 12222 18216
rect 13538 18164 13544 18216
rect 13596 18164 13602 18216
rect 13722 18164 13728 18216
rect 13780 18164 13786 18216
rect 13906 18164 13912 18216
rect 13964 18204 13970 18216
rect 14752 18213 14780 18368
rect 14001 18207 14059 18213
rect 14001 18204 14013 18207
rect 13964 18176 14013 18204
rect 13964 18164 13970 18176
rect 14001 18173 14013 18176
rect 14047 18173 14059 18207
rect 14001 18167 14059 18173
rect 14737 18207 14795 18213
rect 14737 18173 14749 18207
rect 14783 18173 14795 18207
rect 14737 18167 14795 18173
rect 12440 18158 12492 18164
rect 12342 18136 12348 18148
rect 11020 18108 12348 18136
rect 11020 18096 11026 18108
rect 12342 18096 12348 18108
rect 12400 18096 12406 18148
rect 13357 18139 13415 18145
rect 13357 18105 13369 18139
rect 13403 18136 13415 18139
rect 13740 18136 13768 18164
rect 14844 18136 14872 18371
rect 14918 18368 14924 18380
rect 14976 18368 14982 18420
rect 20438 18368 20444 18420
rect 20496 18368 20502 18420
rect 21634 18408 21640 18420
rect 20732 18380 21640 18408
rect 16482 18340 16488 18352
rect 16040 18312 16488 18340
rect 15197 18275 15255 18281
rect 15197 18241 15209 18275
rect 15243 18272 15255 18275
rect 15473 18275 15531 18281
rect 15473 18272 15485 18275
rect 15243 18244 15485 18272
rect 15243 18241 15255 18244
rect 15197 18235 15255 18241
rect 15473 18241 15485 18244
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 15930 18164 15936 18216
rect 15988 18204 15994 18216
rect 16040 18213 16068 18312
rect 16482 18300 16488 18312
rect 16540 18340 16546 18352
rect 16540 18312 16988 18340
rect 16540 18300 16546 18312
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18241 16175 18275
rect 16117 18235 16175 18241
rect 16025 18207 16083 18213
rect 16025 18204 16037 18207
rect 15988 18176 16037 18204
rect 15988 18164 15994 18176
rect 16025 18173 16037 18176
rect 16071 18173 16083 18207
rect 16132 18204 16160 18235
rect 16390 18204 16396 18216
rect 16132 18176 16396 18204
rect 16025 18167 16083 18173
rect 16390 18164 16396 18176
rect 16448 18164 16454 18216
rect 16960 18213 16988 18312
rect 20456 18272 20484 18368
rect 20732 18352 20760 18380
rect 21634 18368 21640 18380
rect 21692 18368 21698 18420
rect 21818 18368 21824 18420
rect 21876 18417 21882 18420
rect 21876 18411 21925 18417
rect 21876 18377 21879 18411
rect 21913 18377 21925 18411
rect 21876 18371 21925 18377
rect 22005 18411 22063 18417
rect 22005 18377 22017 18411
rect 22051 18408 22063 18411
rect 22094 18408 22100 18420
rect 22051 18380 22100 18408
rect 22051 18377 22063 18380
rect 22005 18371 22063 18377
rect 21876 18368 21882 18371
rect 22094 18368 22100 18380
rect 22152 18368 22158 18420
rect 20714 18340 20720 18352
rect 20640 18312 20720 18340
rect 20640 18281 20668 18312
rect 20714 18300 20720 18312
rect 20772 18300 20778 18352
rect 21085 18343 21143 18349
rect 21085 18309 21097 18343
rect 21131 18340 21143 18343
rect 22646 18340 22652 18352
rect 21131 18312 22652 18340
rect 21131 18309 21143 18312
rect 21085 18303 21143 18309
rect 22646 18300 22652 18312
rect 22704 18300 22710 18352
rect 20533 18275 20591 18281
rect 20533 18272 20545 18275
rect 20456 18244 20545 18272
rect 20533 18241 20545 18244
rect 20579 18241 20591 18275
rect 20533 18235 20591 18241
rect 20625 18275 20683 18281
rect 20625 18241 20637 18275
rect 20671 18241 20683 18275
rect 20993 18275 21051 18281
rect 20993 18272 21005 18275
rect 20625 18235 20683 18241
rect 20732 18244 21005 18272
rect 20732 18216 20760 18244
rect 20993 18241 21005 18244
rect 21039 18241 21051 18275
rect 20993 18235 21051 18241
rect 22094 18232 22100 18284
rect 22152 18232 22158 18284
rect 22373 18275 22431 18281
rect 22373 18272 22385 18275
rect 22204 18244 22385 18272
rect 16945 18207 17003 18213
rect 16945 18173 16957 18207
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 17310 18164 17316 18216
rect 17368 18164 17374 18216
rect 20714 18164 20720 18216
rect 20772 18164 20778 18216
rect 20806 18164 20812 18216
rect 20864 18164 20870 18216
rect 21450 18164 21456 18216
rect 21508 18164 21514 18216
rect 22204 18213 22232 18244
rect 22373 18241 22385 18244
rect 22419 18241 22431 18275
rect 22373 18235 22431 18241
rect 21729 18207 21787 18213
rect 21729 18173 21741 18207
rect 21775 18173 21787 18207
rect 21729 18167 21787 18173
rect 22189 18207 22247 18213
rect 22189 18173 22201 18207
rect 22235 18173 22247 18207
rect 22189 18167 22247 18173
rect 22281 18207 22339 18213
rect 22281 18173 22293 18207
rect 22327 18173 22339 18207
rect 22465 18207 22523 18213
rect 22465 18204 22477 18207
rect 22281 18167 22339 18173
rect 22388 18176 22477 18204
rect 16850 18136 16856 18148
rect 13403 18108 13768 18136
rect 14108 18108 14872 18136
rect 16040 18108 16856 18136
rect 13403 18105 13415 18108
rect 13357 18099 13415 18105
rect 4890 18068 4896 18080
rect 4448 18040 4896 18068
rect 4890 18028 4896 18040
rect 4948 18028 4954 18080
rect 7374 18028 7380 18080
rect 7432 18028 7438 18080
rect 8386 18028 8392 18080
rect 8444 18028 8450 18080
rect 10689 18071 10747 18077
rect 10689 18037 10701 18071
rect 10735 18068 10747 18071
rect 14108 18068 14136 18108
rect 10735 18040 14136 18068
rect 14185 18071 14243 18077
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 14185 18037 14197 18071
rect 14231 18068 14243 18071
rect 14550 18068 14556 18080
rect 14231 18040 14556 18068
rect 14231 18037 14243 18040
rect 14185 18031 14243 18037
rect 14550 18028 14556 18040
rect 14608 18028 14614 18080
rect 16040 18077 16068 18108
rect 16850 18096 16856 18108
rect 16908 18096 16914 18148
rect 21358 18096 21364 18148
rect 21416 18136 21422 18148
rect 21416 18108 21496 18136
rect 21416 18096 21422 18108
rect 16025 18071 16083 18077
rect 16025 18037 16037 18071
rect 16071 18037 16083 18071
rect 16025 18031 16083 18037
rect 16301 18071 16359 18077
rect 16301 18037 16313 18071
rect 16347 18068 16359 18071
rect 16574 18068 16580 18080
rect 16347 18040 16580 18068
rect 16347 18037 16359 18040
rect 16301 18031 16359 18037
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 20346 18028 20352 18080
rect 20404 18028 20410 18080
rect 21468 18077 21496 18108
rect 21744 18080 21772 18167
rect 21818 18096 21824 18148
rect 21876 18136 21882 18148
rect 22296 18136 22324 18167
rect 21876 18108 22324 18136
rect 21876 18096 21882 18108
rect 21453 18071 21511 18077
rect 21453 18037 21465 18071
rect 21499 18037 21511 18071
rect 21453 18031 21511 18037
rect 21634 18028 21640 18080
rect 21692 18028 21698 18080
rect 21726 18028 21732 18080
rect 21784 18068 21790 18080
rect 22388 18068 22416 18176
rect 22465 18173 22477 18176
rect 22511 18173 22523 18207
rect 22465 18167 22523 18173
rect 21784 18040 22416 18068
rect 21784 18028 21790 18040
rect 552 17978 23368 18000
rect 552 17926 19022 17978
rect 19074 17926 19086 17978
rect 19138 17926 19150 17978
rect 19202 17926 19214 17978
rect 19266 17926 19278 17978
rect 19330 17926 23368 17978
rect 552 17904 23368 17926
rect 5169 17867 5227 17873
rect 5169 17833 5181 17867
rect 5215 17864 5227 17867
rect 5994 17864 6000 17876
rect 5215 17836 6000 17864
rect 5215 17833 5227 17836
rect 5169 17827 5227 17833
rect 5994 17824 6000 17836
rect 6052 17824 6058 17876
rect 8294 17824 8300 17876
rect 8352 17824 8358 17876
rect 13357 17867 13415 17873
rect 13357 17833 13369 17867
rect 13403 17833 13415 17867
rect 13357 17827 13415 17833
rect 13541 17867 13599 17873
rect 13541 17833 13553 17867
rect 13587 17864 13599 17867
rect 13722 17864 13728 17876
rect 13587 17836 13728 17864
rect 13587 17833 13599 17836
rect 13541 17827 13599 17833
rect 6917 17799 6975 17805
rect 6917 17765 6929 17799
rect 6963 17796 6975 17799
rect 8941 17799 8999 17805
rect 6963 17768 8800 17796
rect 6963 17765 6975 17768
rect 6917 17759 6975 17765
rect 4801 17731 4859 17737
rect 4801 17697 4813 17731
rect 4847 17728 4859 17731
rect 4890 17728 4896 17740
rect 4847 17700 4896 17728
rect 4847 17697 4859 17700
rect 4801 17691 4859 17697
rect 4890 17688 4896 17700
rect 4948 17688 4954 17740
rect 5810 17688 5816 17740
rect 5868 17728 5874 17740
rect 5905 17731 5963 17737
rect 5905 17728 5917 17731
rect 5868 17700 5917 17728
rect 5868 17688 5874 17700
rect 5905 17697 5917 17700
rect 5951 17697 5963 17731
rect 5905 17691 5963 17697
rect 6454 17688 6460 17740
rect 6512 17688 6518 17740
rect 7374 17688 7380 17740
rect 7432 17728 7438 17740
rect 7929 17731 7987 17737
rect 7929 17728 7941 17731
rect 7432 17700 7941 17728
rect 7432 17688 7438 17700
rect 7929 17697 7941 17700
rect 7975 17697 7987 17731
rect 7929 17691 7987 17697
rect 8113 17731 8171 17737
rect 8113 17697 8125 17731
rect 8159 17697 8171 17731
rect 8113 17691 8171 17697
rect 4706 17620 4712 17672
rect 4764 17620 4770 17672
rect 8128 17592 8156 17691
rect 8202 17688 8208 17740
rect 8260 17688 8266 17740
rect 8772 17737 8800 17768
rect 8941 17765 8953 17799
rect 8987 17796 8999 17799
rect 13372 17796 13400 17827
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 13814 17824 13820 17876
rect 13872 17864 13878 17876
rect 15930 17864 15936 17876
rect 13872 17836 15936 17864
rect 13872 17824 13878 17836
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 18782 17824 18788 17876
rect 18840 17824 18846 17876
rect 19610 17824 19616 17876
rect 19668 17873 19674 17876
rect 19668 17827 19677 17873
rect 20441 17867 20499 17873
rect 20441 17833 20453 17867
rect 20487 17864 20499 17867
rect 20806 17864 20812 17876
rect 20487 17836 20812 17864
rect 20487 17833 20499 17836
rect 20441 17827 20499 17833
rect 19668 17824 19674 17827
rect 20806 17824 20812 17836
rect 20864 17824 20870 17876
rect 21361 17867 21419 17873
rect 21361 17833 21373 17867
rect 21407 17864 21419 17867
rect 21450 17864 21456 17876
rect 21407 17836 21456 17864
rect 21407 17833 21419 17836
rect 21361 17827 21419 17833
rect 21450 17824 21456 17836
rect 21508 17824 21514 17876
rect 21637 17867 21695 17873
rect 21637 17833 21649 17867
rect 21683 17864 21695 17867
rect 21818 17864 21824 17876
rect 21683 17836 21824 17864
rect 21683 17833 21695 17836
rect 21637 17827 21695 17833
rect 21818 17824 21824 17836
rect 21876 17824 21882 17876
rect 8987 17768 11836 17796
rect 13372 17768 13676 17796
rect 8987 17765 8999 17768
rect 8941 17759 8999 17765
rect 8757 17731 8815 17737
rect 8757 17697 8769 17731
rect 8803 17728 8815 17731
rect 9125 17731 9183 17737
rect 9125 17728 9137 17731
rect 8803 17700 9137 17728
rect 8803 17697 8815 17700
rect 8757 17691 8815 17697
rect 9125 17697 9137 17700
rect 9171 17697 9183 17731
rect 9125 17691 9183 17697
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 9456 17700 9505 17728
rect 9456 17688 9462 17700
rect 9493 17697 9505 17700
rect 9539 17728 9551 17731
rect 9858 17728 9864 17740
rect 9539 17700 9864 17728
rect 9539 17697 9551 17700
rect 9493 17691 9551 17697
rect 9858 17688 9864 17700
rect 9916 17688 9922 17740
rect 10870 17728 10876 17740
rect 9968 17700 10876 17728
rect 8665 17663 8723 17669
rect 8665 17629 8677 17663
rect 8711 17660 8723 17663
rect 9968 17660 9996 17700
rect 10870 17688 10876 17700
rect 10928 17688 10934 17740
rect 11072 17669 11100 17768
rect 11149 17731 11207 17737
rect 11149 17697 11161 17731
rect 11195 17728 11207 17731
rect 11238 17728 11244 17740
rect 11195 17700 11244 17728
rect 11195 17697 11207 17700
rect 11149 17691 11207 17697
rect 11238 17688 11244 17700
rect 11296 17728 11302 17740
rect 11808 17737 11836 17768
rect 11609 17731 11667 17737
rect 11609 17728 11621 17731
rect 11296 17700 11621 17728
rect 11296 17688 11302 17700
rect 11609 17697 11621 17700
rect 11655 17697 11667 17731
rect 11609 17691 11667 17697
rect 11793 17731 11851 17737
rect 11793 17697 11805 17731
rect 11839 17697 11851 17731
rect 13538 17728 13544 17740
rect 13499 17700 13544 17728
rect 11793 17691 11851 17697
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 8711 17632 9996 17660
rect 10045 17663 10103 17669
rect 8711 17629 8723 17632
rect 8665 17623 8723 17629
rect 10045 17629 10057 17663
rect 10091 17629 10103 17663
rect 10045 17623 10103 17629
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 8680 17592 8708 17623
rect 8128 17564 8708 17592
rect 10060 17536 10088 17623
rect 13556 17592 13584 17688
rect 13648 17660 13676 17768
rect 13740 17728 13768 17824
rect 14277 17731 14335 17737
rect 13740 17700 14228 17728
rect 13906 17660 13912 17672
rect 13648 17632 13912 17660
rect 13906 17620 13912 17632
rect 13964 17620 13970 17672
rect 14001 17663 14059 17669
rect 14001 17629 14013 17663
rect 14047 17660 14059 17663
rect 14090 17660 14096 17672
rect 14047 17632 14096 17660
rect 14047 17629 14059 17632
rect 14001 17623 14059 17629
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14200 17669 14228 17700
rect 14277 17697 14289 17731
rect 14323 17697 14335 17731
rect 15948 17728 15976 17824
rect 18800 17796 18828 17824
rect 19334 17796 19340 17808
rect 18708 17768 18828 17796
rect 18984 17768 19340 17796
rect 18708 17737 18736 17768
rect 18984 17737 19012 17768
rect 19334 17756 19340 17768
rect 19392 17756 19398 17808
rect 19426 17756 19432 17808
rect 19484 17796 19490 17808
rect 19521 17799 19579 17805
rect 19521 17796 19533 17799
rect 19484 17768 19533 17796
rect 19484 17756 19490 17768
rect 19521 17765 19533 17768
rect 19567 17765 19579 17799
rect 21726 17796 21732 17808
rect 19521 17759 19579 17765
rect 20272 17768 21732 17796
rect 20272 17740 20300 17768
rect 16485 17731 16543 17737
rect 16485 17728 16497 17731
rect 15948 17700 16497 17728
rect 14277 17691 14335 17697
rect 16485 17697 16497 17700
rect 16531 17697 16543 17731
rect 16485 17691 16543 17697
rect 18693 17731 18751 17737
rect 18693 17697 18705 17731
rect 18739 17697 18751 17731
rect 18693 17691 18751 17697
rect 18785 17731 18843 17737
rect 18785 17697 18797 17731
rect 18831 17697 18843 17731
rect 18785 17691 18843 17697
rect 18969 17731 19027 17737
rect 18969 17697 18981 17731
rect 19015 17697 19027 17731
rect 18969 17691 19027 17697
rect 14185 17663 14243 17669
rect 14185 17629 14197 17663
rect 14231 17629 14243 17663
rect 14185 17623 14243 17629
rect 14292 17592 14320 17691
rect 16390 17620 16396 17672
rect 16448 17620 16454 17672
rect 18601 17663 18659 17669
rect 18601 17629 18613 17663
rect 18647 17660 18659 17663
rect 18800 17660 18828 17691
rect 19058 17688 19064 17740
rect 19116 17688 19122 17740
rect 19150 17688 19156 17740
rect 19208 17688 19214 17740
rect 19705 17731 19763 17737
rect 19705 17697 19717 17731
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 19720 17660 19748 17691
rect 18647 17632 19748 17660
rect 18647 17629 18659 17632
rect 18601 17623 18659 17629
rect 13556 17564 14320 17592
rect 14645 17595 14703 17601
rect 14645 17561 14657 17595
rect 14691 17592 14703 17595
rect 15102 17592 15108 17604
rect 14691 17564 15108 17592
rect 14691 17561 14703 17564
rect 14645 17555 14703 17561
rect 15102 17552 15108 17564
rect 15160 17552 15166 17604
rect 18966 17552 18972 17604
rect 19024 17592 19030 17604
rect 19812 17592 19840 17691
rect 20254 17688 20260 17740
rect 20312 17688 20318 17740
rect 20809 17731 20867 17737
rect 20809 17697 20821 17731
rect 20855 17728 20867 17731
rect 20990 17728 20996 17740
rect 20855 17700 20996 17728
rect 20855 17697 20867 17700
rect 20809 17691 20867 17697
rect 20990 17688 20996 17700
rect 21048 17688 21054 17740
rect 21284 17737 21312 17768
rect 21726 17756 21732 17768
rect 21784 17756 21790 17808
rect 22278 17756 22284 17808
rect 22336 17796 22342 17808
rect 22750 17799 22808 17805
rect 22750 17796 22762 17799
rect 22336 17768 22762 17796
rect 22336 17756 22342 17768
rect 22750 17765 22762 17768
rect 22796 17765 22808 17799
rect 22750 17759 22808 17765
rect 21269 17731 21327 17737
rect 21269 17697 21281 17731
rect 21315 17697 21327 17731
rect 21269 17691 21327 17697
rect 21358 17688 21364 17740
rect 21416 17688 21422 17740
rect 21453 17731 21511 17737
rect 21453 17697 21465 17731
rect 21499 17728 21511 17731
rect 21542 17728 21548 17740
rect 21499 17700 21548 17728
rect 21499 17697 21511 17700
rect 21453 17691 21511 17697
rect 21542 17688 21548 17700
rect 21600 17688 21606 17740
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17660 20131 17663
rect 20530 17660 20536 17672
rect 20119 17632 20536 17660
rect 20119 17629 20131 17632
rect 20073 17623 20131 17629
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 20625 17663 20683 17669
rect 20625 17629 20637 17663
rect 20671 17629 20683 17663
rect 20625 17623 20683 17629
rect 19024 17564 19840 17592
rect 20640 17592 20668 17623
rect 20714 17620 20720 17672
rect 20772 17620 20778 17672
rect 20901 17663 20959 17669
rect 20901 17629 20913 17663
rect 20947 17660 20959 17663
rect 21376 17660 21404 17688
rect 20947 17632 21404 17660
rect 20947 17629 20959 17632
rect 20901 17623 20959 17629
rect 23014 17620 23020 17672
rect 23072 17620 23078 17672
rect 21358 17592 21364 17604
rect 20640 17564 21364 17592
rect 19024 17552 19030 17564
rect 21358 17552 21364 17564
rect 21416 17552 21422 17604
rect 7742 17484 7748 17536
rect 7800 17484 7806 17536
rect 10042 17484 10048 17536
rect 10100 17484 10106 17536
rect 11514 17484 11520 17536
rect 11572 17484 11578 17536
rect 11974 17484 11980 17536
rect 12032 17484 12038 17536
rect 13909 17527 13967 17533
rect 13909 17493 13921 17527
rect 13955 17524 13967 17527
rect 14274 17524 14280 17536
rect 13955 17496 14280 17524
rect 13955 17493 13967 17496
rect 13909 17487 13967 17493
rect 14274 17484 14280 17496
rect 14332 17484 14338 17536
rect 16206 17484 16212 17536
rect 16264 17484 16270 17536
rect 18230 17484 18236 17536
rect 18288 17524 18294 17536
rect 19150 17524 19156 17536
rect 18288 17496 19156 17524
rect 18288 17484 18294 17496
rect 19150 17484 19156 17496
rect 19208 17484 19214 17536
rect 19429 17527 19487 17533
rect 19429 17493 19441 17527
rect 19475 17524 19487 17527
rect 20622 17524 20628 17536
rect 19475 17496 20628 17524
rect 19475 17493 19487 17496
rect 19429 17487 19487 17493
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 21082 17484 21088 17536
rect 21140 17484 21146 17536
rect 552 17434 23368 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 23368 17434
rect 552 17360 23368 17382
rect 7742 17280 7748 17332
rect 7800 17280 7806 17332
rect 11974 17280 11980 17332
rect 12032 17280 12038 17332
rect 12158 17280 12164 17332
rect 12216 17280 12222 17332
rect 14274 17280 14280 17332
rect 14332 17320 14338 17332
rect 14553 17323 14611 17329
rect 14553 17320 14565 17323
rect 14332 17292 14565 17320
rect 14332 17280 14338 17292
rect 14553 17289 14565 17292
rect 14599 17289 14611 17323
rect 14553 17283 14611 17289
rect 16206 17280 16212 17332
rect 16264 17280 16270 17332
rect 16485 17323 16543 17329
rect 16485 17289 16497 17323
rect 16531 17320 16543 17323
rect 16666 17320 16672 17332
rect 16531 17292 16672 17320
rect 16531 17289 16543 17292
rect 16485 17283 16543 17289
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 18782 17280 18788 17332
rect 18840 17280 18846 17332
rect 18966 17280 18972 17332
rect 19024 17280 19030 17332
rect 19058 17280 19064 17332
rect 19116 17280 19122 17332
rect 21082 17280 21088 17332
rect 21140 17280 21146 17332
rect 21358 17280 21364 17332
rect 21416 17320 21422 17332
rect 22649 17323 22707 17329
rect 22649 17320 22661 17323
rect 21416 17292 22661 17320
rect 21416 17280 21422 17292
rect 22649 17289 22661 17292
rect 22695 17289 22707 17323
rect 22649 17283 22707 17289
rect 7760 17252 7788 17280
rect 7760 17224 9628 17252
rect 8202 17144 8208 17196
rect 8260 17184 8266 17196
rect 8757 17187 8815 17193
rect 8757 17184 8769 17187
rect 8260 17156 8769 17184
rect 8260 17144 8266 17156
rect 8757 17153 8769 17156
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 8849 17119 8907 17125
rect 8849 17085 8861 17119
rect 8895 17116 8907 17119
rect 9398 17116 9404 17128
rect 8895 17088 9404 17116
rect 8895 17085 8907 17088
rect 8849 17079 8907 17085
rect 9398 17076 9404 17088
rect 9456 17076 9462 17128
rect 9600 17048 9628 17224
rect 9677 17187 9735 17193
rect 9677 17153 9689 17187
rect 9723 17184 9735 17187
rect 10042 17184 10048 17196
rect 9723 17156 10048 17184
rect 9723 17153 9735 17156
rect 9677 17147 9735 17153
rect 10042 17144 10048 17156
rect 10100 17184 10106 17196
rect 11425 17187 11483 17193
rect 10100 17156 10824 17184
rect 10100 17144 10106 17156
rect 10796 17125 10824 17156
rect 11425 17153 11437 17187
rect 11471 17184 11483 17187
rect 11514 17184 11520 17196
rect 11471 17156 11520 17184
rect 11471 17153 11483 17156
rect 11425 17147 11483 17153
rect 11514 17144 11520 17156
rect 11572 17184 11578 17196
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 11572 17156 11805 17184
rect 11572 17144 11578 17156
rect 11793 17153 11805 17156
rect 11839 17153 11851 17187
rect 11992 17184 12020 17280
rect 12176 17252 12204 17280
rect 16224 17252 16252 17280
rect 17405 17255 17463 17261
rect 17405 17252 17417 17255
rect 12176 17224 14688 17252
rect 12345 17187 12403 17193
rect 12345 17184 12357 17187
rect 11992 17156 12357 17184
rect 11793 17147 11851 17153
rect 12345 17153 12357 17156
rect 12391 17153 12403 17187
rect 12345 17147 12403 17153
rect 13909 17187 13967 17193
rect 13909 17153 13921 17187
rect 13955 17184 13967 17187
rect 14274 17184 14280 17196
rect 13955 17156 14280 17184
rect 13955 17153 13967 17156
rect 13909 17147 13967 17153
rect 14274 17144 14280 17156
rect 14332 17144 14338 17196
rect 10597 17119 10655 17125
rect 10597 17116 10609 17119
rect 10166 17102 10609 17116
rect 10152 17088 10609 17102
rect 10152 17048 10180 17088
rect 10597 17085 10609 17088
rect 10643 17085 10655 17119
rect 10597 17079 10655 17085
rect 10781 17119 10839 17125
rect 10781 17085 10793 17119
rect 10827 17085 10839 17119
rect 10781 17079 10839 17085
rect 11333 17119 11391 17125
rect 11333 17085 11345 17119
rect 11379 17116 11391 17119
rect 11977 17119 12035 17125
rect 11977 17116 11989 17119
rect 11379 17088 11989 17116
rect 11379 17085 11391 17088
rect 11333 17079 11391 17085
rect 9600 17020 10180 17048
rect 10505 17051 10563 17057
rect 10505 17017 10517 17051
rect 10551 17048 10563 17051
rect 11146 17048 11152 17060
rect 10551 17020 11152 17048
rect 10551 17017 10563 17020
rect 10505 17011 10563 17017
rect 11146 17008 11152 17020
rect 11204 17008 11210 17060
rect 11440 16992 11468 17088
rect 11977 17085 11989 17088
rect 12023 17116 12035 17119
rect 13814 17116 13820 17128
rect 12023 17088 13820 17116
rect 12023 17085 12035 17088
rect 11977 17079 12035 17085
rect 13814 17076 13820 17088
rect 13872 17076 13878 17128
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17116 14059 17119
rect 14090 17116 14096 17128
rect 14047 17088 14096 17116
rect 14047 17085 14059 17088
rect 14001 17079 14059 17085
rect 14090 17076 14096 17088
rect 14148 17116 14154 17128
rect 14461 17119 14519 17125
rect 14461 17116 14473 17119
rect 14148 17088 14473 17116
rect 14148 17076 14154 17088
rect 14461 17085 14473 17088
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 14550 17076 14556 17128
rect 14608 17076 14614 17128
rect 14660 17116 14688 17224
rect 16132 17224 16252 17252
rect 16684 17224 17417 17252
rect 14734 17144 14740 17196
rect 14792 17144 14798 17196
rect 16025 17187 16083 17193
rect 16025 17184 16037 17187
rect 15672 17156 16037 17184
rect 15672 17125 15700 17156
rect 16025 17153 16037 17156
rect 16071 17153 16083 17187
rect 16025 17147 16083 17153
rect 16132 17125 16160 17224
rect 16684 17125 16712 17224
rect 17405 17221 17417 17224
rect 17451 17221 17463 17255
rect 17405 17215 17463 17221
rect 17494 17212 17500 17264
rect 17552 17252 17558 17264
rect 18800 17252 18828 17280
rect 17552 17224 17908 17252
rect 18800 17224 18920 17252
rect 17552 17212 17558 17224
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 17328 17156 17785 17184
rect 15657 17119 15715 17125
rect 15657 17116 15669 17119
rect 14660 17088 15669 17116
rect 15657 17085 15669 17088
rect 15703 17085 15715 17119
rect 15657 17079 15715 17085
rect 15841 17119 15899 17125
rect 15841 17085 15853 17119
rect 15887 17116 15899 17119
rect 16117 17119 16175 17125
rect 16117 17116 16129 17119
rect 15887 17088 16129 17116
rect 15887 17085 15899 17088
rect 15841 17079 15899 17085
rect 16117 17085 16129 17088
rect 16163 17085 16175 17119
rect 16117 17079 16175 17085
rect 16669 17119 16727 17125
rect 16669 17085 16681 17119
rect 16715 17085 16727 17119
rect 16669 17079 16727 17085
rect 16762 17119 16820 17125
rect 16762 17085 16774 17119
rect 16808 17085 16820 17119
rect 16762 17079 16820 17085
rect 17175 17119 17233 17125
rect 17175 17085 17187 17119
rect 17221 17116 17233 17119
rect 17328 17116 17356 17156
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 17773 17147 17831 17153
rect 17221 17088 17356 17116
rect 17221 17085 17233 17088
rect 17175 17079 17233 17085
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 13170 17048 13176 17060
rect 12584 17020 13176 17048
rect 12584 17008 12590 17020
rect 13170 17008 13176 17020
rect 13228 17008 13234 17060
rect 13262 17008 13268 17060
rect 13320 17048 13326 17060
rect 14182 17048 14188 17060
rect 13320 17020 14188 17048
rect 13320 17008 13326 17020
rect 14182 17008 14188 17020
rect 14240 17008 14246 17060
rect 14568 17048 14596 17076
rect 15930 17048 15936 17060
rect 14568 17020 15936 17048
rect 15930 17008 15936 17020
rect 15988 17048 15994 17060
rect 16776 17048 16804 17079
rect 17402 17076 17408 17128
rect 17460 17076 17466 17128
rect 17880 17125 17908 17224
rect 18892 17125 18920 17224
rect 18984 17193 19012 17280
rect 18969 17187 19027 17193
rect 18969 17153 18981 17187
rect 19015 17153 19027 17187
rect 18969 17147 19027 17153
rect 17589 17119 17647 17125
rect 17589 17085 17601 17119
rect 17635 17116 17647 17119
rect 17681 17119 17739 17125
rect 17681 17116 17693 17119
rect 17635 17088 17693 17116
rect 17635 17085 17647 17088
rect 17589 17079 17647 17085
rect 17681 17085 17693 17088
rect 17727 17085 17739 17119
rect 17681 17079 17739 17085
rect 17865 17119 17923 17125
rect 17865 17085 17877 17119
rect 17911 17085 17923 17119
rect 17865 17079 17923 17085
rect 18877 17119 18935 17125
rect 18877 17085 18889 17119
rect 18923 17085 18935 17119
rect 18877 17079 18935 17085
rect 15988 17020 16804 17048
rect 15988 17008 15994 17020
rect 16942 17008 16948 17060
rect 17000 17008 17006 17060
rect 17037 17051 17095 17057
rect 17037 17017 17049 17051
rect 17083 17017 17095 17051
rect 17604 17048 17632 17079
rect 17037 17011 17095 17017
rect 17144 17020 17632 17048
rect 18141 17051 18199 17057
rect 9214 16940 9220 16992
rect 9272 16940 9278 16992
rect 10778 16940 10784 16992
rect 10836 16940 10842 16992
rect 11422 16940 11428 16992
rect 11480 16940 11486 16992
rect 11698 16940 11704 16992
rect 11756 16940 11762 16992
rect 12158 16940 12164 16992
rect 12216 16980 12222 16992
rect 12253 16983 12311 16989
rect 12253 16980 12265 16983
rect 12216 16952 12265 16980
rect 12216 16940 12222 16952
rect 12253 16949 12265 16952
rect 12299 16949 12311 16983
rect 12253 16943 12311 16949
rect 14366 16940 14372 16992
rect 14424 16940 14430 16992
rect 14737 16983 14795 16989
rect 14737 16949 14749 16983
rect 14783 16980 14795 16983
rect 15010 16980 15016 16992
rect 14783 16952 15016 16980
rect 14783 16949 14795 16952
rect 14737 16943 14795 16949
rect 15010 16940 15016 16952
rect 15068 16940 15074 16992
rect 15749 16983 15807 16989
rect 15749 16949 15761 16983
rect 15795 16980 15807 16983
rect 16758 16980 16764 16992
rect 15795 16952 16764 16980
rect 15795 16949 15807 16952
rect 15749 16943 15807 16949
rect 16758 16940 16764 16952
rect 16816 16980 16822 16992
rect 17052 16980 17080 17011
rect 17144 16992 17172 17020
rect 18141 17017 18153 17051
rect 18187 17017 18199 17051
rect 18141 17011 18199 17017
rect 16816 16952 17080 16980
rect 16816 16940 16822 16952
rect 17126 16940 17132 16992
rect 17184 16940 17190 16992
rect 17313 16983 17371 16989
rect 17313 16949 17325 16983
rect 17359 16980 17371 16983
rect 18156 16980 18184 17011
rect 18230 17008 18236 17060
rect 18288 17048 18294 17060
rect 18325 17051 18383 17057
rect 18325 17048 18337 17051
rect 18288 17020 18337 17048
rect 18288 17008 18294 17020
rect 18325 17017 18337 17020
rect 18371 17017 18383 17051
rect 18325 17011 18383 17017
rect 18509 17051 18567 17057
rect 18509 17017 18521 17051
rect 18555 17048 18567 17051
rect 18984 17048 19012 17147
rect 18555 17020 19012 17048
rect 18555 17017 18567 17020
rect 18509 17011 18567 17017
rect 19076 16980 19104 17280
rect 21100 17184 21128 17280
rect 22186 17212 22192 17264
rect 22244 17252 22250 17264
rect 22557 17255 22615 17261
rect 22557 17252 22569 17255
rect 22244 17224 22569 17252
rect 22244 17212 22250 17224
rect 22557 17221 22569 17224
rect 22603 17252 22615 17255
rect 22603 17224 23060 17252
rect 22603 17221 22615 17224
rect 22557 17215 22615 17221
rect 23032 17193 23060 17224
rect 23017 17187 23075 17193
rect 21100 17156 21312 17184
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17116 19763 17119
rect 19794 17116 19800 17128
rect 19751 17088 19800 17116
rect 19751 17085 19763 17088
rect 19705 17079 19763 17085
rect 19794 17076 19800 17088
rect 19852 17076 19858 17128
rect 19972 17119 20030 17125
rect 19972 17085 19984 17119
rect 20018 17116 20030 17119
rect 20346 17116 20352 17128
rect 20018 17088 20352 17116
rect 20018 17085 20030 17088
rect 19972 17079 20030 17085
rect 20346 17076 20352 17088
rect 20404 17076 20410 17128
rect 20530 17076 20536 17128
rect 20588 17076 20594 17128
rect 21174 17076 21180 17128
rect 21232 17076 21238 17128
rect 21284 17116 21312 17156
rect 23017 17153 23029 17187
rect 23063 17153 23075 17187
rect 23017 17147 23075 17153
rect 21433 17119 21491 17125
rect 21433 17116 21445 17119
rect 21284 17088 21445 17116
rect 21433 17085 21445 17088
rect 21479 17085 21491 17119
rect 21433 17079 21491 17085
rect 21726 17076 21732 17128
rect 21784 17116 21790 17128
rect 22833 17119 22891 17125
rect 22833 17116 22845 17119
rect 21784 17088 22845 17116
rect 21784 17076 21790 17088
rect 22833 17085 22845 17088
rect 22879 17085 22891 17119
rect 22833 17079 22891 17085
rect 17359 16952 19104 16980
rect 19245 16983 19303 16989
rect 17359 16949 17371 16952
rect 17313 16943 17371 16949
rect 19245 16949 19257 16983
rect 19291 16980 19303 16983
rect 20070 16980 20076 16992
rect 19291 16952 20076 16980
rect 19291 16949 19303 16952
rect 19245 16943 19303 16949
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 20548 16980 20576 17076
rect 21085 16983 21143 16989
rect 21085 16980 21097 16983
rect 20548 16952 21097 16980
rect 21085 16949 21097 16952
rect 21131 16949 21143 16983
rect 21085 16943 21143 16949
rect 552 16890 23368 16912
rect 552 16838 19022 16890
rect 19074 16838 19086 16890
rect 19138 16838 19150 16890
rect 19202 16838 19214 16890
rect 19266 16838 19278 16890
rect 19330 16838 23368 16890
rect 552 16816 23368 16838
rect 7006 16736 7012 16788
rect 7064 16736 7070 16788
rect 10229 16779 10287 16785
rect 10229 16745 10241 16779
rect 10275 16745 10287 16779
rect 10229 16739 10287 16745
rect 6089 16711 6147 16717
rect 6089 16677 6101 16711
rect 6135 16708 6147 16711
rect 6135 16680 6684 16708
rect 6135 16677 6147 16680
rect 6089 16671 6147 16677
rect 5997 16643 6055 16649
rect 5997 16609 6009 16643
rect 6043 16640 6055 16643
rect 6273 16643 6331 16649
rect 6043 16612 6224 16640
rect 6043 16609 6055 16612
rect 5997 16603 6055 16609
rect 6196 16584 6224 16612
rect 6273 16609 6285 16643
rect 6319 16640 6331 16643
rect 6454 16640 6460 16652
rect 6319 16612 6460 16640
rect 6319 16609 6331 16612
rect 6273 16603 6331 16609
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16609 6607 16643
rect 6549 16603 6607 16609
rect 6178 16532 6184 16584
rect 6236 16532 6242 16584
rect 6564 16448 6592 16603
rect 6656 16572 6684 16680
rect 6733 16643 6791 16649
rect 6733 16609 6745 16643
rect 6779 16640 6791 16643
rect 6822 16640 6828 16652
rect 6779 16612 6828 16640
rect 6779 16609 6791 16612
rect 6733 16603 6791 16609
rect 6822 16600 6828 16612
rect 6880 16640 6886 16652
rect 7024 16640 7052 16736
rect 9214 16668 9220 16720
rect 9272 16708 9278 16720
rect 9769 16711 9827 16717
rect 9769 16708 9781 16711
rect 9272 16680 9781 16708
rect 9272 16668 9278 16680
rect 9769 16677 9781 16680
rect 9815 16677 9827 16711
rect 9769 16671 9827 16677
rect 6880 16612 7052 16640
rect 10244 16640 10272 16739
rect 10778 16736 10784 16788
rect 10836 16776 10842 16788
rect 10836 16748 11008 16776
rect 10836 16736 10842 16748
rect 10980 16717 11008 16748
rect 11514 16736 11520 16788
rect 11572 16736 11578 16788
rect 12526 16736 12532 16788
rect 12584 16736 12590 16788
rect 13262 16776 13268 16788
rect 12636 16748 13268 16776
rect 10965 16711 11023 16717
rect 10965 16677 10977 16711
rect 11011 16677 11023 16711
rect 12636 16708 12664 16748
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 14734 16736 14740 16788
rect 14792 16736 14798 16788
rect 16850 16736 16856 16788
rect 16908 16776 16914 16788
rect 17402 16776 17408 16788
rect 16908 16748 17408 16776
rect 16908 16736 16914 16748
rect 17402 16736 17408 16748
rect 17460 16736 17466 16788
rect 19426 16736 19432 16788
rect 19484 16736 19490 16788
rect 22646 16736 22652 16788
rect 22704 16736 22710 16788
rect 19444 16708 19472 16736
rect 10965 16671 11023 16677
rect 12406 16680 12664 16708
rect 18892 16680 19472 16708
rect 21536 16711 21594 16717
rect 11054 16640 11060 16652
rect 10244 16612 11060 16640
rect 6880 16600 6886 16612
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 11146 16600 11152 16652
rect 11204 16600 11210 16652
rect 11422 16600 11428 16652
rect 11480 16640 11486 16652
rect 11517 16643 11575 16649
rect 11517 16640 11529 16643
rect 11480 16612 11529 16640
rect 11480 16600 11486 16612
rect 11517 16609 11529 16612
rect 11563 16609 11575 16643
rect 11517 16603 11575 16609
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16640 12127 16643
rect 12406 16640 12434 16680
rect 12618 16649 12624 16652
rect 12115 16612 12434 16640
rect 12588 16643 12624 16649
rect 12115 16609 12127 16612
rect 12069 16603 12127 16609
rect 12588 16609 12600 16643
rect 12676 16640 12682 16652
rect 13449 16643 13507 16649
rect 13449 16640 13461 16643
rect 12676 16612 13461 16640
rect 12588 16603 12624 16609
rect 12618 16600 12624 16603
rect 12676 16600 12682 16612
rect 13449 16609 13461 16612
rect 13495 16640 13507 16643
rect 14001 16643 14059 16649
rect 14001 16640 14013 16643
rect 13495 16612 14013 16640
rect 13495 16609 13507 16612
rect 13449 16603 13507 16609
rect 14001 16609 14013 16612
rect 14047 16609 14059 16643
rect 14185 16643 14243 16649
rect 14185 16640 14197 16643
rect 14001 16603 14059 16609
rect 14108 16612 14197 16640
rect 11164 16572 11192 16600
rect 11609 16575 11667 16581
rect 11609 16572 11621 16575
rect 6656 16544 6960 16572
rect 11164 16544 11621 16572
rect 6932 16448 6960 16544
rect 11609 16541 11621 16544
rect 11655 16541 11667 16575
rect 11609 16535 11667 16541
rect 11882 16532 11888 16584
rect 11940 16532 11946 16584
rect 12897 16575 12955 16581
rect 12897 16541 12909 16575
rect 12943 16572 12955 16575
rect 13078 16572 13084 16584
rect 12943 16544 13084 16572
rect 12943 16541 12955 16544
rect 12897 16535 12955 16541
rect 13078 16532 13084 16544
rect 13136 16532 13142 16584
rect 13170 16532 13176 16584
rect 13228 16572 13234 16584
rect 13357 16575 13415 16581
rect 13357 16572 13369 16575
rect 13228 16544 13369 16572
rect 13228 16532 13234 16544
rect 13357 16541 13369 16544
rect 13403 16572 13415 16575
rect 14108 16572 14136 16612
rect 14185 16609 14197 16612
rect 14231 16609 14243 16643
rect 14461 16643 14519 16649
rect 14461 16640 14473 16643
rect 14185 16603 14243 16609
rect 14292 16612 14473 16640
rect 13403 16544 14136 16572
rect 13403 16541 13415 16544
rect 13357 16535 13415 16541
rect 9490 16464 9496 16516
rect 9548 16504 9554 16516
rect 10045 16507 10103 16513
rect 10045 16504 10057 16507
rect 9548 16476 10057 16504
rect 9548 16464 9554 16476
rect 10045 16473 10057 16476
rect 10091 16473 10103 16507
rect 10045 16467 10103 16473
rect 6457 16439 6515 16445
rect 6457 16405 6469 16439
rect 6503 16436 6515 16439
rect 6546 16436 6552 16448
rect 6503 16408 6552 16436
rect 6503 16405 6515 16408
rect 6457 16399 6515 16405
rect 6546 16396 6552 16408
rect 6604 16396 6610 16448
rect 6638 16396 6644 16448
rect 6696 16396 6702 16448
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 11900 16436 11928 16532
rect 12713 16507 12771 16513
rect 12713 16473 12725 16507
rect 12759 16504 12771 16507
rect 14292 16504 14320 16612
rect 14461 16609 14473 16612
rect 14507 16609 14519 16643
rect 14461 16603 14519 16609
rect 15197 16643 15255 16649
rect 15197 16609 15209 16643
rect 15243 16640 15255 16643
rect 15654 16640 15660 16652
rect 15243 16612 15660 16640
rect 15243 16609 15255 16612
rect 15197 16603 15255 16609
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 16669 16643 16727 16649
rect 16669 16640 16681 16643
rect 16632 16612 16681 16640
rect 16632 16600 16638 16612
rect 16669 16609 16681 16612
rect 16715 16640 16727 16643
rect 17126 16640 17132 16652
rect 16715 16612 17132 16640
rect 16715 16609 16727 16612
rect 16669 16603 16727 16609
rect 17126 16600 17132 16612
rect 17184 16600 17190 16652
rect 18892 16649 18920 16680
rect 21536 16677 21548 16711
rect 21582 16708 21594 16711
rect 21634 16708 21640 16720
rect 21582 16680 21640 16708
rect 21582 16677 21594 16680
rect 21536 16671 21594 16677
rect 21634 16668 21640 16680
rect 21692 16668 21698 16720
rect 17313 16643 17371 16649
rect 17313 16609 17325 16643
rect 17359 16609 17371 16643
rect 17313 16603 17371 16609
rect 18877 16643 18935 16649
rect 18877 16609 18889 16643
rect 18923 16609 18935 16643
rect 19610 16640 19616 16652
rect 18877 16603 18935 16609
rect 18984 16612 19616 16640
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 16761 16575 16819 16581
rect 14424 16544 15056 16572
rect 14424 16532 14430 16544
rect 12759 16476 14320 16504
rect 12759 16473 12771 16476
rect 12713 16467 12771 16473
rect 6972 16408 11928 16436
rect 6972 16396 6978 16408
rect 12158 16396 12164 16448
rect 12216 16396 12222 16448
rect 13906 16396 13912 16448
rect 13964 16436 13970 16448
rect 14384 16436 14412 16532
rect 13964 16408 14412 16436
rect 13964 16396 13970 16408
rect 14642 16396 14648 16448
rect 14700 16396 14706 16448
rect 14918 16396 14924 16448
rect 14976 16436 14982 16448
rect 15028 16445 15056 16544
rect 16761 16541 16773 16575
rect 16807 16572 16819 16575
rect 16850 16572 16856 16584
rect 16807 16544 16856 16572
rect 16807 16541 16819 16544
rect 16761 16535 16819 16541
rect 16850 16532 16856 16544
rect 16908 16532 16914 16584
rect 17034 16532 17040 16584
rect 17092 16572 17098 16584
rect 17328 16572 17356 16603
rect 18984 16581 19012 16612
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 19794 16600 19800 16652
rect 19852 16640 19858 16652
rect 23014 16640 23020 16652
rect 19852 16612 23020 16640
rect 19852 16600 19858 16612
rect 23014 16600 23020 16612
rect 23072 16600 23078 16652
rect 17092 16544 17356 16572
rect 17497 16575 17555 16581
rect 17092 16532 17098 16544
rect 17497 16541 17509 16575
rect 17543 16541 17555 16575
rect 17497 16535 17555 16541
rect 18969 16575 19027 16581
rect 18969 16541 18981 16575
rect 19015 16541 19027 16575
rect 18969 16535 19027 16541
rect 16666 16464 16672 16516
rect 16724 16504 16730 16516
rect 17512 16504 17540 16535
rect 21174 16532 21180 16584
rect 21232 16572 21238 16584
rect 21269 16575 21327 16581
rect 21269 16572 21281 16575
rect 21232 16544 21281 16572
rect 21232 16532 21238 16544
rect 21269 16541 21281 16544
rect 21315 16541 21327 16575
rect 21269 16535 21327 16541
rect 16724 16476 17540 16504
rect 16724 16464 16730 16476
rect 15013 16439 15071 16445
rect 15013 16436 15025 16439
rect 14976 16408 15025 16436
rect 14976 16396 14982 16408
rect 15013 16405 15025 16408
rect 15059 16405 15071 16439
rect 15013 16399 15071 16405
rect 16574 16396 16580 16448
rect 16632 16436 16638 16448
rect 16942 16436 16948 16448
rect 16632 16408 16948 16436
rect 16632 16396 16638 16408
rect 16942 16396 16948 16408
rect 17000 16436 17006 16448
rect 17129 16439 17187 16445
rect 17129 16436 17141 16439
rect 17000 16408 17141 16436
rect 17000 16396 17006 16408
rect 17129 16405 17141 16408
rect 17175 16405 17187 16439
rect 17129 16399 17187 16405
rect 18874 16396 18880 16448
rect 18932 16436 18938 16448
rect 19153 16439 19211 16445
rect 19153 16436 19165 16439
rect 18932 16408 19165 16436
rect 18932 16396 18938 16408
rect 19153 16405 19165 16408
rect 19199 16405 19211 16439
rect 19153 16399 19211 16405
rect 552 16346 23368 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 23368 16346
rect 552 16272 23368 16294
rect 6178 16232 6184 16244
rect 4816 16204 6184 16232
rect 4816 16037 4844 16204
rect 6178 16192 6184 16204
rect 6236 16192 6242 16244
rect 9490 16192 9496 16244
rect 9548 16232 9554 16244
rect 10045 16235 10103 16241
rect 10045 16232 10057 16235
rect 9548 16204 10057 16232
rect 9548 16192 9554 16204
rect 5077 16167 5135 16173
rect 5077 16133 5089 16167
rect 5123 16133 5135 16167
rect 5077 16127 5135 16133
rect 5092 16096 5120 16127
rect 6454 16124 6460 16176
rect 6512 16164 6518 16176
rect 6512 16136 7420 16164
rect 6512 16124 6518 16136
rect 5092 16068 5764 16096
rect 4801 16031 4859 16037
rect 4801 15997 4813 16031
rect 4847 15997 4859 16031
rect 4801 15991 4859 15997
rect 5074 15988 5080 16040
rect 5132 16028 5138 16040
rect 5736 16037 5764 16068
rect 6362 16056 6368 16108
rect 6420 16096 6426 16108
rect 6914 16096 6920 16108
rect 6420 16068 6920 16096
rect 6420 16056 6426 16068
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 5353 16031 5411 16037
rect 5353 16028 5365 16031
rect 5132 16000 5365 16028
rect 5132 15988 5138 16000
rect 5353 15997 5365 16000
rect 5399 15997 5411 16031
rect 5353 15991 5411 15997
rect 5445 16031 5503 16037
rect 5445 15997 5457 16031
rect 5491 16028 5503 16031
rect 5721 16031 5779 16037
rect 5491 16000 5672 16028
rect 5491 15997 5503 16000
rect 5445 15991 5503 15997
rect 4893 15963 4951 15969
rect 4893 15929 4905 15963
rect 4939 15960 4951 15963
rect 4939 15932 5488 15960
rect 4939 15929 4951 15932
rect 4893 15923 4951 15929
rect 5460 15904 5488 15932
rect 5534 15920 5540 15972
rect 5592 15920 5598 15972
rect 5644 15960 5672 16000
rect 5721 15997 5733 16031
rect 5767 15997 5779 16031
rect 5721 15991 5779 15997
rect 5902 15988 5908 16040
rect 5960 16028 5966 16040
rect 5997 16031 6055 16037
rect 5997 16028 6009 16031
rect 5960 16000 6009 16028
rect 5960 15988 5966 16000
rect 5997 15997 6009 16000
rect 6043 15997 6055 16031
rect 5997 15991 6055 15997
rect 6454 15988 6460 16040
rect 6512 15988 6518 16040
rect 6638 15988 6644 16040
rect 6696 16028 6702 16040
rect 6733 16031 6791 16037
rect 6733 16028 6745 16031
rect 6696 16000 6745 16028
rect 6696 15988 6702 16000
rect 6733 15997 6745 16000
rect 6779 15997 6791 16031
rect 6733 15991 6791 15997
rect 5644 15932 6040 15960
rect 6012 15904 6040 15932
rect 6086 15920 6092 15972
rect 6144 15920 6150 15972
rect 6932 15969 6960 16056
rect 7024 16037 7052 16136
rect 7285 16099 7343 16105
rect 7285 16065 7297 16099
rect 7331 16065 7343 16099
rect 7285 16059 7343 16065
rect 7009 16031 7067 16037
rect 7009 15997 7021 16031
rect 7055 15997 7067 16031
rect 7009 15991 7067 15997
rect 6181 15963 6239 15969
rect 6181 15929 6193 15963
rect 6227 15929 6239 15963
rect 6181 15923 6239 15929
rect 6299 15963 6357 15969
rect 6299 15929 6311 15963
rect 6345 15960 6357 15963
rect 6917 15963 6975 15969
rect 6345 15932 6776 15960
rect 6345 15929 6357 15932
rect 6299 15923 6357 15929
rect 5166 15852 5172 15904
rect 5224 15852 5230 15904
rect 5442 15852 5448 15904
rect 5500 15852 5506 15904
rect 5626 15852 5632 15904
rect 5684 15892 5690 15904
rect 5813 15895 5871 15901
rect 5813 15892 5825 15895
rect 5684 15864 5825 15892
rect 5684 15852 5690 15864
rect 5813 15861 5825 15864
rect 5859 15861 5871 15895
rect 5813 15855 5871 15861
rect 5994 15852 6000 15904
rect 6052 15852 6058 15904
rect 6196 15892 6224 15923
rect 6748 15904 6776 15932
rect 6917 15929 6929 15963
rect 6963 15929 6975 15963
rect 6917 15923 6975 15929
rect 7300 15904 7328 16059
rect 7392 15960 7420 16136
rect 7558 16056 7564 16108
rect 7616 16096 7622 16108
rect 8018 16096 8024 16108
rect 7616 16068 8024 16096
rect 7616 16056 7622 16068
rect 8018 16056 8024 16068
rect 8076 16056 8082 16108
rect 9600 16105 9628 16204
rect 10045 16201 10057 16204
rect 10091 16201 10103 16235
rect 15102 16232 15108 16244
rect 10045 16195 10103 16201
rect 14108 16204 15108 16232
rect 9585 16099 9643 16105
rect 9585 16065 9597 16099
rect 9631 16065 9643 16099
rect 9585 16059 9643 16065
rect 11146 16056 11152 16108
rect 11204 16056 11210 16108
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 16028 7711 16031
rect 7834 16028 7840 16040
rect 7699 16000 7840 16028
rect 7699 15997 7711 16000
rect 7653 15991 7711 15997
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 9214 15988 9220 16040
rect 9272 16028 9278 16040
rect 9493 16031 9551 16037
rect 9493 16028 9505 16031
rect 9272 16000 9505 16028
rect 9272 15988 9278 16000
rect 9493 15997 9505 16000
rect 9539 16028 9551 16031
rect 9953 16031 10011 16037
rect 9953 16028 9965 16031
rect 9539 16000 9965 16028
rect 9539 15997 9551 16000
rect 9493 15991 9551 15997
rect 9953 15997 9965 16000
rect 9999 15997 10011 16031
rect 9953 15991 10011 15997
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 16028 11115 16031
rect 11422 16028 11428 16040
rect 11103 16000 11428 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 11422 15988 11428 16000
rect 11480 15988 11486 16040
rect 13906 15988 13912 16040
rect 13964 15988 13970 16040
rect 14108 16037 14136 16204
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 21913 16235 21971 16241
rect 21913 16201 21925 16235
rect 21959 16232 21971 16235
rect 22094 16232 22100 16244
rect 21959 16204 22100 16232
rect 21959 16201 21971 16204
rect 21913 16195 21971 16201
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 22925 16235 22983 16241
rect 22925 16201 22937 16235
rect 22971 16232 22983 16235
rect 23014 16232 23020 16244
rect 22971 16204 23020 16232
rect 22971 16201 22983 16204
rect 22925 16195 22983 16201
rect 14461 16167 14519 16173
rect 14461 16133 14473 16167
rect 14507 16164 14519 16167
rect 14642 16164 14648 16176
rect 14507 16136 14648 16164
rect 14507 16133 14519 16136
rect 14461 16127 14519 16133
rect 14642 16124 14648 16136
rect 14700 16124 14706 16176
rect 16574 16164 16580 16176
rect 14844 16136 16580 16164
rect 14093 16031 14151 16037
rect 14093 15997 14105 16031
rect 14139 15997 14151 16031
rect 14093 15991 14151 15997
rect 14366 15988 14372 16040
rect 14424 15988 14430 16040
rect 14550 15988 14556 16040
rect 14608 15988 14614 16040
rect 14844 16037 14872 16136
rect 16574 16124 16580 16136
rect 16632 16124 16638 16176
rect 16761 16167 16819 16173
rect 16761 16133 16773 16167
rect 16807 16133 16819 16167
rect 22940 16164 22968 16195
rect 23014 16192 23020 16204
rect 23072 16192 23078 16244
rect 16761 16127 16819 16133
rect 22296 16136 22968 16164
rect 15010 16056 15016 16108
rect 15068 16056 15074 16108
rect 16776 16096 16804 16127
rect 16945 16099 17003 16105
rect 16945 16096 16957 16099
rect 16776 16068 16957 16096
rect 16945 16065 16957 16068
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 14645 16031 14703 16037
rect 14645 15997 14657 16031
rect 14691 15997 14703 16031
rect 14645 15991 14703 15997
rect 14829 16031 14887 16037
rect 14829 15997 14841 16031
rect 14875 15997 14887 16031
rect 14829 15991 14887 15997
rect 14001 15963 14059 15969
rect 7392 15932 7696 15960
rect 7668 15904 7696 15932
rect 14001 15929 14013 15963
rect 14047 15960 14059 15963
rect 14660 15960 14688 15991
rect 15102 15988 15108 16040
rect 15160 15988 15166 16040
rect 15565 16031 15623 16037
rect 15565 16028 15577 16031
rect 15212 16000 15577 16028
rect 15212 15960 15240 16000
rect 15565 15997 15577 16000
rect 15611 15997 15623 16031
rect 15565 15991 15623 15997
rect 15841 16031 15899 16037
rect 15841 15997 15853 16031
rect 15887 16028 15899 16031
rect 15930 16028 15936 16040
rect 15887 16000 15936 16028
rect 15887 15997 15899 16000
rect 15841 15991 15899 15997
rect 15930 15988 15936 16000
rect 15988 15988 15994 16040
rect 16025 16031 16083 16037
rect 16025 15997 16037 16031
rect 16071 16028 16083 16031
rect 16390 16028 16396 16040
rect 16071 16000 16396 16028
rect 16071 15997 16083 16000
rect 16025 15991 16083 15997
rect 16390 15988 16396 16000
rect 16448 16028 16454 16040
rect 16485 16031 16543 16037
rect 16485 16028 16497 16031
rect 16448 16000 16497 16028
rect 16448 15988 16454 16000
rect 16485 15997 16497 16000
rect 16531 15997 16543 16031
rect 16485 15991 16543 15997
rect 16577 16031 16635 16037
rect 16577 15997 16589 16031
rect 16623 16028 16635 16031
rect 16666 16028 16672 16040
rect 16623 16000 16672 16028
rect 16623 15997 16635 16000
rect 16577 15991 16635 15997
rect 16666 15988 16672 16000
rect 16724 15988 16730 16040
rect 16758 15988 16764 16040
rect 16816 15988 16822 16040
rect 17034 15988 17040 16040
rect 17092 15988 17098 16040
rect 22296 16037 22324 16136
rect 22370 16056 22376 16108
rect 22428 16096 22434 16108
rect 22465 16099 22523 16105
rect 22465 16096 22477 16099
rect 22428 16068 22477 16096
rect 22428 16056 22434 16068
rect 22465 16065 22477 16068
rect 22511 16065 22523 16099
rect 22465 16059 22523 16065
rect 22281 16031 22339 16037
rect 22281 15997 22293 16031
rect 22327 15997 22339 16031
rect 22281 15991 22339 15997
rect 22741 16031 22799 16037
rect 22741 15997 22753 16031
rect 22787 16028 22799 16031
rect 22830 16028 22836 16040
rect 22787 16000 22836 16028
rect 22787 15997 22799 16000
rect 22741 15991 22799 15997
rect 22830 15988 22836 16000
rect 22888 15988 22894 16040
rect 18230 15960 18236 15972
rect 14047 15932 15240 15960
rect 15304 15932 18236 15960
rect 14047 15929 14059 15932
rect 14001 15923 14059 15929
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 6196 15864 6561 15892
rect 6549 15861 6561 15864
rect 6595 15861 6607 15895
rect 6549 15855 6607 15861
rect 6730 15852 6736 15904
rect 6788 15852 6794 15904
rect 7282 15852 7288 15904
rect 7340 15852 7346 15904
rect 7650 15852 7656 15904
rect 7708 15852 7714 15904
rect 9858 15852 9864 15904
rect 9916 15852 9922 15904
rect 10410 15852 10416 15904
rect 10468 15852 10474 15904
rect 11790 15852 11796 15904
rect 11848 15852 11854 15904
rect 14185 15895 14243 15901
rect 14185 15861 14197 15895
rect 14231 15892 14243 15895
rect 15304 15892 15332 15932
rect 18230 15920 18236 15932
rect 18288 15920 18294 15972
rect 22002 15920 22008 15972
rect 22060 15960 22066 15972
rect 22373 15963 22431 15969
rect 22373 15960 22385 15963
rect 22060 15932 22385 15960
rect 22060 15920 22066 15932
rect 22373 15929 22385 15932
rect 22419 15929 22431 15963
rect 22373 15923 22431 15929
rect 14231 15864 15332 15892
rect 14231 15861 14243 15864
rect 14185 15855 14243 15861
rect 15470 15852 15476 15904
rect 15528 15852 15534 15904
rect 15654 15852 15660 15904
rect 15712 15852 15718 15904
rect 17402 15852 17408 15904
rect 17460 15852 17466 15904
rect 552 15802 23368 15824
rect 552 15750 19022 15802
rect 19074 15750 19086 15802
rect 19138 15750 19150 15802
rect 19202 15750 19214 15802
rect 19266 15750 19278 15802
rect 19330 15750 23368 15802
rect 552 15728 23368 15750
rect 5166 15648 5172 15700
rect 5224 15648 5230 15700
rect 5534 15648 5540 15700
rect 5592 15688 5598 15700
rect 5813 15691 5871 15697
rect 5813 15688 5825 15691
rect 5592 15660 5825 15688
rect 5592 15648 5598 15660
rect 5813 15657 5825 15660
rect 5859 15657 5871 15691
rect 5813 15651 5871 15657
rect 5902 15648 5908 15700
rect 5960 15648 5966 15700
rect 6086 15648 6092 15700
rect 6144 15688 6150 15700
rect 6273 15691 6331 15697
rect 6273 15688 6285 15691
rect 6144 15660 6285 15688
rect 6144 15648 6150 15660
rect 6273 15657 6285 15660
rect 6319 15657 6331 15691
rect 6825 15691 6883 15697
rect 6825 15688 6837 15691
rect 6273 15651 6331 15657
rect 6472 15660 6837 15688
rect 4516 15623 4574 15629
rect 4516 15589 4528 15623
rect 4562 15620 4574 15623
rect 5184 15620 5212 15648
rect 4562 15592 5212 15620
rect 5920 15620 5948 15648
rect 6472 15620 6500 15660
rect 6825 15657 6837 15660
rect 6871 15657 6883 15691
rect 6825 15651 6883 15657
rect 9858 15648 9864 15700
rect 9916 15648 9922 15700
rect 10410 15648 10416 15700
rect 10468 15648 10474 15700
rect 14366 15688 14372 15700
rect 13464 15660 14372 15688
rect 5920 15592 6500 15620
rect 4562 15589 4574 15592
rect 4516 15583 4574 15589
rect 6546 15580 6552 15632
rect 6604 15620 6610 15632
rect 6641 15623 6699 15629
rect 6641 15620 6653 15623
rect 6604 15592 6653 15620
rect 6604 15580 6610 15592
rect 6641 15589 6653 15592
rect 6687 15589 6699 15623
rect 7282 15620 7288 15632
rect 6641 15583 6699 15589
rect 7208 15592 7288 15620
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 5997 15555 6055 15561
rect 5997 15552 6009 15555
rect 5592 15524 6009 15552
rect 5592 15512 5598 15524
rect 5997 15521 6009 15524
rect 6043 15521 6055 15555
rect 5997 15515 6055 15521
rect 4249 15487 4307 15493
rect 4249 15453 4261 15487
rect 4295 15453 4307 15487
rect 6012 15484 6040 15515
rect 6178 15512 6184 15564
rect 6236 15512 6242 15564
rect 6362 15512 6368 15564
rect 6420 15512 6426 15564
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15521 6515 15555
rect 6457 15515 6515 15521
rect 6380 15484 6408 15512
rect 6012 15456 6408 15484
rect 6472 15484 6500 15515
rect 6730 15512 6736 15564
rect 6788 15512 6794 15564
rect 6822 15512 6828 15564
rect 6880 15512 6886 15564
rect 7208 15561 7236 15592
rect 7282 15580 7288 15592
rect 7340 15620 7346 15632
rect 7340 15592 8524 15620
rect 7340 15580 7346 15592
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15521 6975 15555
rect 6917 15515 6975 15521
rect 7009 15555 7067 15561
rect 7009 15521 7021 15555
rect 7055 15521 7067 15555
rect 7009 15515 7067 15521
rect 7193 15555 7251 15561
rect 7193 15521 7205 15555
rect 7239 15521 7251 15555
rect 7193 15515 7251 15521
rect 7469 15555 7527 15561
rect 7469 15521 7481 15555
rect 7515 15552 7527 15555
rect 7515 15524 7972 15552
rect 7515 15521 7527 15524
rect 7469 15515 7527 15521
rect 6840 15484 6868 15512
rect 6472 15456 6868 15484
rect 4249 15447 4307 15453
rect 4264 15348 4292 15447
rect 6932 15416 6960 15515
rect 7024 15484 7052 15515
rect 7484 15484 7512 15515
rect 7024 15456 7512 15484
rect 7650 15444 7656 15496
rect 7708 15444 7714 15496
rect 7834 15444 7840 15496
rect 7892 15444 7898 15496
rect 7944 15484 7972 15524
rect 8018 15512 8024 15564
rect 8076 15512 8082 15564
rect 8496 15561 8524 15592
rect 8481 15555 8539 15561
rect 8481 15521 8493 15555
rect 8527 15521 8539 15555
rect 8481 15515 8539 15521
rect 8665 15487 8723 15493
rect 8665 15484 8677 15487
rect 7944 15456 8677 15484
rect 8665 15453 8677 15456
rect 8711 15453 8723 15487
rect 9876 15484 9904 15648
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15521 10195 15555
rect 10428 15552 10456 15648
rect 13464 15564 13492 15660
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 16390 15648 16396 15700
rect 16448 15648 16454 15700
rect 18874 15648 18880 15700
rect 18932 15688 18938 15700
rect 19061 15691 19119 15697
rect 19061 15688 19073 15691
rect 18932 15660 19073 15688
rect 18932 15648 18938 15660
rect 19061 15657 19073 15660
rect 19107 15657 19119 15691
rect 19061 15651 19119 15657
rect 20070 15648 20076 15700
rect 20128 15648 20134 15700
rect 16408 15620 16436 15648
rect 17313 15623 17371 15629
rect 17313 15620 17325 15623
rect 13556 15592 14688 15620
rect 11241 15555 11299 15561
rect 11241 15552 11253 15555
rect 10428 15524 11253 15552
rect 10137 15515 10195 15521
rect 11241 15521 11253 15524
rect 11287 15521 11299 15555
rect 12986 15552 12992 15564
rect 11241 15515 11299 15521
rect 12406 15524 12992 15552
rect 10045 15487 10103 15493
rect 10045 15484 10057 15487
rect 9876 15456 10057 15484
rect 8665 15447 8723 15453
rect 10045 15453 10057 15456
rect 10091 15453 10103 15487
rect 10152 15484 10180 15515
rect 10962 15484 10968 15496
rect 10152 15456 10968 15484
rect 10045 15447 10103 15453
rect 7852 15416 7880 15444
rect 8680 15416 8708 15447
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11054 15444 11060 15496
rect 11112 15444 11118 15496
rect 12406 15416 12434 15524
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 13170 15512 13176 15564
rect 13228 15512 13234 15564
rect 13446 15512 13452 15564
rect 13504 15512 13510 15564
rect 13556 15561 13584 15592
rect 14660 15564 14688 15592
rect 16408 15592 17325 15620
rect 13541 15555 13599 15561
rect 13541 15521 13553 15555
rect 13587 15521 13599 15555
rect 13541 15515 13599 15521
rect 13725 15555 13783 15561
rect 13725 15521 13737 15555
rect 13771 15521 13783 15555
rect 13725 15515 13783 15521
rect 13817 15555 13875 15561
rect 13817 15521 13829 15555
rect 13863 15552 13875 15555
rect 14550 15552 14556 15564
rect 13863 15524 14556 15552
rect 13863 15521 13875 15524
rect 13817 15515 13875 15521
rect 12526 15444 12532 15496
rect 12584 15484 12590 15496
rect 13740 15484 13768 15515
rect 12584 15456 13768 15484
rect 12584 15444 12590 15456
rect 6932 15388 7328 15416
rect 7852 15388 8432 15416
rect 8680 15388 12434 15416
rect 13357 15419 13415 15425
rect 4522 15348 4528 15360
rect 4264 15320 4528 15348
rect 4522 15308 4528 15320
rect 4580 15308 4586 15360
rect 5629 15351 5687 15357
rect 5629 15317 5641 15351
rect 5675 15348 5687 15351
rect 5994 15348 6000 15360
rect 5675 15320 6000 15348
rect 5675 15317 5687 15320
rect 5629 15311 5687 15317
rect 5994 15308 6000 15320
rect 6052 15308 6058 15360
rect 7190 15308 7196 15360
rect 7248 15308 7254 15360
rect 7300 15357 7328 15388
rect 7285 15351 7343 15357
rect 7285 15317 7297 15351
rect 7331 15348 7343 15351
rect 7742 15348 7748 15360
rect 7331 15320 7748 15348
rect 7331 15317 7343 15320
rect 7285 15311 7343 15317
rect 7742 15308 7748 15320
rect 7800 15308 7806 15360
rect 8202 15308 8208 15360
rect 8260 15308 8266 15360
rect 8294 15308 8300 15360
rect 8352 15308 8358 15360
rect 8404 15348 8432 15388
rect 13357 15385 13369 15419
rect 13403 15416 13415 15419
rect 13832 15416 13860 15515
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 14642 15512 14648 15564
rect 14700 15512 14706 15564
rect 14829 15555 14887 15561
rect 14829 15521 14841 15555
rect 14875 15552 14887 15555
rect 14918 15552 14924 15564
rect 14875 15524 14924 15552
rect 14875 15521 14887 15524
rect 14829 15515 14887 15521
rect 14918 15512 14924 15524
rect 14976 15512 14982 15564
rect 16408 15561 16436 15592
rect 17313 15589 17325 15592
rect 17359 15589 17371 15623
rect 17313 15583 17371 15589
rect 21174 15580 21180 15632
rect 21232 15620 21238 15632
rect 22830 15620 22836 15632
rect 21232 15592 22836 15620
rect 21232 15580 21238 15592
rect 22830 15580 22836 15592
rect 22888 15580 22894 15632
rect 16393 15555 16451 15561
rect 16393 15521 16405 15555
rect 16439 15521 16451 15555
rect 16393 15515 16451 15521
rect 16577 15555 16635 15561
rect 16577 15521 16589 15555
rect 16623 15552 16635 15555
rect 16666 15552 16672 15564
rect 16623 15524 16672 15552
rect 16623 15521 16635 15524
rect 16577 15515 16635 15521
rect 16666 15512 16672 15524
rect 16724 15552 16730 15564
rect 17497 15555 17555 15561
rect 17497 15552 17509 15555
rect 16724 15524 17509 15552
rect 16724 15512 16730 15524
rect 17497 15521 17509 15524
rect 17543 15521 17555 15555
rect 17497 15515 17555 15521
rect 18414 15512 18420 15564
rect 18472 15552 18478 15564
rect 19153 15555 19211 15561
rect 19153 15552 19165 15555
rect 18472 15524 19165 15552
rect 18472 15512 18478 15524
rect 19153 15521 19165 15524
rect 19199 15521 19211 15555
rect 19153 15515 19211 15521
rect 19978 15512 19984 15564
rect 20036 15512 20042 15564
rect 14001 15487 14059 15493
rect 14001 15453 14013 15487
rect 14047 15484 14059 15487
rect 14737 15487 14795 15493
rect 14737 15484 14749 15487
rect 14047 15456 14749 15484
rect 14047 15453 14059 15456
rect 14001 15447 14059 15453
rect 14737 15453 14749 15456
rect 14783 15484 14795 15487
rect 15654 15484 15660 15496
rect 14783 15456 15660 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 16485 15487 16543 15493
rect 16485 15453 16497 15487
rect 16531 15484 16543 15487
rect 16853 15487 16911 15493
rect 16853 15484 16865 15487
rect 16531 15456 16865 15484
rect 16531 15453 16543 15456
rect 16485 15447 16543 15453
rect 16853 15453 16865 15456
rect 16899 15453 16911 15487
rect 16853 15447 16911 15453
rect 16945 15487 17003 15493
rect 16945 15453 16957 15487
rect 16991 15453 17003 15487
rect 16945 15447 17003 15453
rect 13403 15388 13860 15416
rect 13403 15385 13415 15388
rect 13357 15379 13415 15385
rect 15194 15376 15200 15428
rect 15252 15376 15258 15428
rect 16960 15416 16988 15447
rect 17034 15444 17040 15496
rect 17092 15444 17098 15496
rect 17129 15487 17187 15493
rect 17129 15453 17141 15487
rect 17175 15484 17187 15487
rect 17770 15484 17776 15496
rect 17175 15456 17776 15484
rect 17175 15453 17187 15456
rect 17129 15447 17187 15453
rect 17770 15444 17776 15456
rect 17828 15444 17834 15496
rect 18969 15487 19027 15493
rect 18969 15453 18981 15487
rect 19015 15484 19027 15487
rect 19426 15484 19432 15496
rect 19015 15456 19432 15484
rect 19015 15453 19027 15456
rect 18969 15447 19027 15453
rect 19426 15444 19432 15456
rect 19484 15484 19490 15496
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 19484 15456 20177 15484
rect 19484 15444 19490 15456
rect 20165 15453 20177 15456
rect 20211 15453 20223 15487
rect 21192 15484 21220 15580
rect 21358 15512 21364 15564
rect 21416 15552 21422 15564
rect 21525 15555 21583 15561
rect 21525 15552 21537 15555
rect 21416 15524 21537 15552
rect 21416 15512 21422 15524
rect 21525 15521 21537 15524
rect 21571 15521 21583 15555
rect 21525 15515 21583 15521
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 21192 15456 21281 15484
rect 20165 15447 20223 15453
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 17681 15419 17739 15425
rect 17681 15416 17693 15419
rect 16960 15388 17693 15416
rect 17681 15385 17693 15388
rect 17727 15385 17739 15419
rect 17681 15379 17739 15385
rect 9030 15348 9036 15360
rect 8404 15320 9036 15348
rect 9030 15308 9036 15320
rect 9088 15308 9094 15360
rect 9858 15308 9864 15360
rect 9916 15308 9922 15360
rect 11422 15308 11428 15360
rect 11480 15308 11486 15360
rect 16574 15308 16580 15360
rect 16632 15348 16638 15360
rect 16669 15351 16727 15357
rect 16669 15348 16681 15351
rect 16632 15320 16681 15348
rect 16632 15308 16638 15320
rect 16669 15317 16681 15320
rect 16715 15317 16727 15351
rect 16669 15311 16727 15317
rect 19518 15308 19524 15360
rect 19576 15308 19582 15360
rect 19610 15308 19616 15360
rect 19668 15308 19674 15360
rect 22002 15308 22008 15360
rect 22060 15348 22066 15360
rect 22649 15351 22707 15357
rect 22649 15348 22661 15351
rect 22060 15320 22661 15348
rect 22060 15308 22066 15320
rect 22649 15317 22661 15320
rect 22695 15317 22707 15351
rect 22649 15311 22707 15317
rect 552 15258 23368 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 23368 15258
rect 552 15184 23368 15206
rect 6273 15147 6331 15153
rect 6273 15113 6285 15147
rect 6319 15144 6331 15147
rect 6454 15144 6460 15156
rect 6319 15116 6460 15144
rect 6319 15113 6331 15116
rect 6273 15107 6331 15113
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 6914 15104 6920 15156
rect 6972 15144 6978 15156
rect 7190 15144 7196 15156
rect 6972 15116 7196 15144
rect 6972 15104 6978 15116
rect 7190 15104 7196 15116
rect 7248 15144 7254 15156
rect 7377 15147 7435 15153
rect 7377 15144 7389 15147
rect 7248 15116 7389 15144
rect 7248 15104 7254 15116
rect 7377 15113 7389 15116
rect 7423 15113 7435 15147
rect 7377 15107 7435 15113
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8573 15147 8631 15153
rect 8573 15144 8585 15147
rect 8352 15116 8585 15144
rect 8352 15104 8358 15116
rect 8573 15113 8585 15116
rect 8619 15113 8631 15147
rect 8573 15107 8631 15113
rect 11422 15104 11428 15156
rect 11480 15144 11486 15156
rect 12069 15147 12127 15153
rect 12069 15144 12081 15147
rect 11480 15116 12081 15144
rect 11480 15104 11486 15116
rect 12069 15113 12081 15116
rect 12115 15113 12127 15147
rect 12069 15107 12127 15113
rect 13173 15147 13231 15153
rect 13173 15113 13185 15147
rect 13219 15144 13231 15147
rect 13446 15144 13452 15156
rect 13219 15116 13452 15144
rect 13219 15113 13231 15116
rect 13173 15107 13231 15113
rect 13446 15104 13452 15116
rect 13504 15104 13510 15156
rect 17770 15104 17776 15156
rect 17828 15104 17834 15156
rect 19610 15144 19616 15156
rect 18340 15116 19616 15144
rect 7742 15036 7748 15088
rect 7800 15076 7806 15088
rect 7800 15048 9260 15076
rect 7800 15036 7806 15048
rect 6638 14968 6644 15020
rect 6696 15008 6702 15020
rect 8386 15008 8392 15020
rect 6696 14980 7236 15008
rect 6696 14968 6702 14980
rect 4522 14900 4528 14952
rect 4580 14940 4586 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4580 14912 4905 14940
rect 4580 14900 4586 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 5160 14943 5218 14949
rect 5160 14909 5172 14943
rect 5206 14940 5218 14943
rect 5626 14940 5632 14952
rect 5206 14912 5632 14940
rect 5206 14909 5218 14912
rect 5160 14903 5218 14909
rect 5626 14900 5632 14912
rect 5684 14900 5690 14952
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 6840 14872 6868 14903
rect 6914 14900 6920 14952
rect 6972 14900 6978 14952
rect 7208 14949 7236 14980
rect 7760 14980 8392 15008
rect 7760 14949 7788 14980
rect 8386 14968 8392 14980
rect 8444 15008 8450 15020
rect 8444 14980 8984 15008
rect 8444 14968 8450 14980
rect 7193 14943 7251 14949
rect 7193 14909 7205 14943
rect 7239 14909 7251 14943
rect 7193 14903 7251 14909
rect 7469 14943 7527 14949
rect 7469 14909 7481 14943
rect 7515 14909 7527 14943
rect 7469 14903 7527 14909
rect 7745 14943 7803 14949
rect 7745 14909 7757 14943
rect 7791 14909 7803 14943
rect 7745 14903 7803 14909
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14909 8079 14943
rect 8021 14903 8079 14909
rect 7484 14872 7512 14903
rect 8036 14872 8064 14903
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 8956 14949 8984 14980
rect 8573 14943 8631 14949
rect 8573 14940 8585 14943
rect 8260 14912 8585 14940
rect 8260 14900 8266 14912
rect 8573 14909 8585 14912
rect 8619 14909 8631 14943
rect 8573 14903 8631 14909
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14909 8999 14943
rect 8941 14903 8999 14909
rect 9030 14900 9036 14952
rect 9088 14900 9094 14952
rect 9232 14949 9260 15048
rect 12158 15036 12164 15088
rect 12216 15076 12222 15088
rect 13906 15076 13912 15088
rect 12216 15048 13912 15076
rect 12216 15036 12222 15048
rect 13906 15036 13912 15048
rect 13964 15076 13970 15088
rect 13964 15048 14136 15076
rect 13964 15036 13970 15048
rect 11609 15011 11667 15017
rect 11609 14977 11621 15011
rect 11655 15008 11667 15011
rect 11698 15008 11704 15020
rect 11655 14980 11704 15008
rect 11655 14977 11667 14980
rect 11609 14971 11667 14977
rect 11698 14968 11704 14980
rect 11756 15008 11762 15020
rect 12066 15008 12072 15020
rect 11756 14980 12072 15008
rect 11756 14968 11762 14980
rect 12066 14968 12072 14980
rect 12124 15008 12130 15020
rect 12124 14980 12296 15008
rect 12124 14968 12130 14980
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 11514 14900 11520 14952
rect 11572 14900 11578 14952
rect 11790 14900 11796 14952
rect 11848 14940 11854 14952
rect 12268 14949 12296 14980
rect 12526 14968 12532 15020
rect 12584 15008 12590 15020
rect 14108 15017 14136 15048
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12584 14980 13001 15008
rect 12584 14968 12590 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 14093 15011 14151 15017
rect 14093 14977 14105 15011
rect 14139 14977 14151 15011
rect 14093 14971 14151 14977
rect 17972 14980 18184 15008
rect 11977 14943 12035 14949
rect 11977 14940 11989 14943
rect 11848 14912 11989 14940
rect 11848 14900 11854 14912
rect 11977 14909 11989 14912
rect 12023 14909 12035 14943
rect 11977 14903 12035 14909
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14909 12311 14943
rect 12253 14903 12311 14909
rect 12345 14943 12403 14949
rect 12345 14909 12357 14943
rect 12391 14909 12403 14943
rect 12345 14903 12403 14909
rect 12897 14943 12955 14949
rect 12897 14909 12909 14943
rect 12943 14940 12955 14943
rect 12943 14912 13584 14940
rect 12943 14909 12955 14912
rect 12897 14903 12955 14909
rect 8294 14872 8300 14884
rect 6840 14844 8300 14872
rect 8294 14832 8300 14844
rect 8352 14832 8358 14884
rect 11532 14872 11560 14900
rect 12360 14872 12388 14903
rect 11532 14844 12388 14872
rect 12802 14832 12808 14884
rect 12860 14832 12866 14884
rect 13078 14832 13084 14884
rect 13136 14872 13142 14884
rect 13173 14875 13231 14881
rect 13173 14872 13185 14875
rect 13136 14844 13185 14872
rect 13136 14832 13142 14844
rect 13173 14841 13185 14844
rect 13219 14841 13231 14875
rect 13173 14835 13231 14841
rect 6730 14764 6736 14816
rect 6788 14804 6794 14816
rect 6917 14807 6975 14813
rect 6917 14804 6929 14807
rect 6788 14776 6929 14804
rect 6788 14764 6794 14776
rect 6917 14773 6929 14776
rect 6963 14773 6975 14807
rect 6917 14767 6975 14773
rect 7006 14764 7012 14816
rect 7064 14764 7070 14816
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 7561 14807 7619 14813
rect 7561 14804 7573 14807
rect 7156 14776 7573 14804
rect 7156 14764 7162 14776
rect 7561 14773 7573 14776
rect 7607 14804 7619 14807
rect 7834 14804 7840 14816
rect 7607 14776 7840 14804
rect 7607 14773 7619 14776
rect 7561 14767 7619 14773
rect 7834 14764 7840 14776
rect 7892 14764 7898 14816
rect 8110 14764 8116 14816
rect 8168 14804 8174 14816
rect 8389 14807 8447 14813
rect 8389 14804 8401 14807
rect 8168 14776 8401 14804
rect 8168 14764 8174 14776
rect 8389 14773 8401 14776
rect 8435 14773 8447 14807
rect 8389 14767 8447 14773
rect 9122 14764 9128 14816
rect 9180 14764 9186 14816
rect 11882 14764 11888 14816
rect 11940 14764 11946 14816
rect 11974 14764 11980 14816
rect 12032 14804 12038 14816
rect 12342 14804 12348 14816
rect 12032 14776 12348 14804
rect 12032 14764 12038 14776
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 13556 14813 13584 14912
rect 14182 14900 14188 14952
rect 14240 14900 14246 14952
rect 16301 14943 16359 14949
rect 16301 14909 16313 14943
rect 16347 14940 16359 14943
rect 16390 14940 16396 14952
rect 16347 14912 16396 14940
rect 16347 14909 16359 14912
rect 16301 14903 16359 14909
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 16574 14949 16580 14952
rect 16568 14940 16580 14949
rect 16535 14912 16580 14940
rect 16568 14903 16580 14912
rect 16574 14900 16580 14903
rect 16632 14900 16638 14952
rect 17972 14949 18000 14980
rect 17957 14943 18015 14949
rect 17957 14909 17969 14943
rect 18003 14909 18015 14943
rect 17957 14903 18015 14909
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14909 18107 14943
rect 18049 14903 18107 14909
rect 13541 14807 13599 14813
rect 13541 14773 13553 14807
rect 13587 14804 13599 14807
rect 13722 14804 13728 14816
rect 13587 14776 13728 14804
rect 13587 14773 13599 14776
rect 13541 14767 13599 14773
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 17678 14764 17684 14816
rect 17736 14804 17742 14816
rect 18064 14804 18092 14903
rect 18156 14872 18184 14980
rect 18340 14949 18368 15116
rect 19610 15104 19616 15116
rect 19668 15104 19674 15156
rect 19978 15104 19984 15156
rect 20036 15144 20042 15156
rect 20073 15147 20131 15153
rect 20073 15144 20085 15147
rect 20036 15116 20085 15144
rect 20036 15104 20042 15116
rect 20073 15113 20085 15116
rect 20119 15113 20131 15147
rect 20073 15107 20131 15113
rect 21358 15104 21364 15156
rect 21416 15104 21422 15156
rect 21453 15011 21511 15017
rect 18432 14980 18828 15008
rect 18325 14943 18383 14949
rect 18325 14909 18337 14943
rect 18371 14909 18383 14943
rect 18325 14903 18383 14909
rect 18432 14872 18460 14980
rect 18690 14900 18696 14952
rect 18748 14900 18754 14952
rect 18800 14940 18828 14980
rect 21453 14977 21465 15011
rect 21499 14977 21511 15011
rect 21453 14971 21511 14977
rect 18800 14912 19472 14940
rect 18938 14875 18996 14881
rect 18938 14872 18950 14875
rect 18156 14844 18460 14872
rect 18524 14844 18950 14872
rect 18524 14813 18552 14844
rect 18938 14841 18950 14844
rect 18984 14841 18996 14875
rect 19444 14872 19472 14912
rect 19518 14900 19524 14952
rect 19576 14940 19582 14952
rect 20349 14943 20407 14949
rect 20349 14940 20361 14943
rect 19576 14912 20361 14940
rect 19576 14900 19582 14912
rect 20349 14909 20361 14912
rect 20395 14909 20407 14943
rect 20349 14903 20407 14909
rect 20714 14900 20720 14952
rect 20772 14940 20778 14952
rect 21177 14943 21235 14949
rect 21177 14940 21189 14943
rect 20772 14912 21189 14940
rect 20772 14900 20778 14912
rect 21177 14909 21189 14912
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 21361 14943 21419 14949
rect 21361 14909 21373 14943
rect 21407 14940 21419 14943
rect 21468 14940 21496 14971
rect 21910 14968 21916 15020
rect 21968 14968 21974 15020
rect 22296 14980 22692 15008
rect 21407 14912 21496 14940
rect 21821 14943 21879 14949
rect 21407 14909 21419 14912
rect 21361 14903 21419 14909
rect 21821 14909 21833 14943
rect 21867 14940 21879 14943
rect 22002 14940 22008 14952
rect 21867 14912 22008 14940
rect 21867 14909 21879 14912
rect 21821 14903 21879 14909
rect 22002 14900 22008 14912
rect 22060 14900 22066 14952
rect 22296 14949 22324 14980
rect 22664 14952 22692 14980
rect 22281 14943 22339 14949
rect 22281 14909 22293 14943
rect 22327 14909 22339 14943
rect 22281 14903 22339 14909
rect 20254 14872 20260 14884
rect 19444 14844 20260 14872
rect 18938 14835 18996 14841
rect 19536 14816 19564 14844
rect 20254 14832 20260 14844
rect 20312 14832 20318 14884
rect 22296 14872 22324 14903
rect 22646 14900 22652 14952
rect 22704 14900 22710 14952
rect 21468 14844 22324 14872
rect 21468 14816 21496 14844
rect 22462 14832 22468 14884
rect 22520 14832 22526 14884
rect 17736 14776 18092 14804
rect 18509 14807 18567 14813
rect 17736 14764 17742 14776
rect 18509 14773 18521 14807
rect 18555 14773 18567 14807
rect 18509 14767 18567 14773
rect 19518 14764 19524 14816
rect 19576 14764 19582 14816
rect 20162 14764 20168 14816
rect 20220 14764 20226 14816
rect 21450 14764 21456 14816
rect 21508 14764 21514 14816
rect 22097 14807 22155 14813
rect 22097 14773 22109 14807
rect 22143 14804 22155 14807
rect 22370 14804 22376 14816
rect 22143 14776 22376 14804
rect 22143 14773 22155 14776
rect 22097 14767 22155 14773
rect 22370 14764 22376 14776
rect 22428 14764 22434 14816
rect 552 14714 23368 14736
rect 552 14662 19022 14714
rect 19074 14662 19086 14714
rect 19138 14662 19150 14714
rect 19202 14662 19214 14714
rect 19266 14662 19278 14714
rect 19330 14662 23368 14714
rect 552 14640 23368 14662
rect 4890 14560 4896 14612
rect 4948 14600 4954 14612
rect 5169 14603 5227 14609
rect 5169 14600 5181 14603
rect 4948 14572 5181 14600
rect 4948 14560 4954 14572
rect 5169 14569 5181 14572
rect 5215 14569 5227 14603
rect 6730 14600 6736 14612
rect 5169 14563 5227 14569
rect 6380 14572 6736 14600
rect 5077 14467 5135 14473
rect 5077 14433 5089 14467
rect 5123 14464 5135 14467
rect 5718 14464 5724 14476
rect 5123 14436 5724 14464
rect 5123 14433 5135 14436
rect 5077 14427 5135 14433
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 6380 14473 6408 14572
rect 6730 14560 6736 14572
rect 6788 14560 6794 14612
rect 7006 14560 7012 14612
rect 7064 14560 7070 14612
rect 7101 14603 7159 14609
rect 7101 14569 7113 14603
rect 7147 14600 7159 14603
rect 9398 14600 9404 14612
rect 7147 14572 9404 14600
rect 7147 14569 7159 14572
rect 7101 14563 7159 14569
rect 9398 14560 9404 14572
rect 9456 14600 9462 14612
rect 9861 14603 9919 14609
rect 9861 14600 9873 14603
rect 9456 14572 9873 14600
rect 9456 14560 9462 14572
rect 9861 14569 9873 14572
rect 9907 14569 9919 14603
rect 9861 14563 9919 14569
rect 10781 14603 10839 14609
rect 10781 14569 10793 14603
rect 10827 14569 10839 14603
rect 11974 14600 11980 14612
rect 10781 14563 10839 14569
rect 11900 14572 11980 14600
rect 7024 14532 7052 14560
rect 6564 14504 7052 14532
rect 6564 14473 6592 14504
rect 7834 14492 7840 14544
rect 7892 14532 7898 14544
rect 8389 14535 8447 14541
rect 8389 14532 8401 14535
rect 7892 14504 8401 14532
rect 7892 14492 7898 14504
rect 8389 14501 8401 14504
rect 8435 14501 8447 14535
rect 9876 14532 9904 14563
rect 10229 14535 10287 14541
rect 10229 14532 10241 14535
rect 9876 14504 10241 14532
rect 8389 14495 8447 14501
rect 10229 14501 10241 14504
rect 10275 14501 10287 14535
rect 10796 14532 10824 14563
rect 11900 14532 11928 14572
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 12066 14560 12072 14612
rect 12124 14560 12130 14612
rect 12802 14600 12808 14612
rect 12268 14572 12808 14600
rect 10796 14504 11928 14532
rect 10229 14495 10287 14501
rect 6365 14467 6423 14473
rect 6365 14433 6377 14467
rect 6411 14433 6423 14467
rect 6365 14427 6423 14433
rect 6549 14467 6607 14473
rect 6549 14433 6561 14467
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 6638 14424 6644 14476
rect 6696 14424 6702 14476
rect 6730 14424 6736 14476
rect 6788 14424 6794 14476
rect 6917 14467 6975 14473
rect 6917 14433 6929 14467
rect 6963 14464 6975 14467
rect 7098 14464 7104 14476
rect 6963 14436 7104 14464
rect 6963 14433 6975 14436
rect 6917 14427 6975 14433
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 7190 14424 7196 14476
rect 7248 14424 7254 14476
rect 7374 14430 7380 14482
rect 7432 14430 7438 14482
rect 7466 14424 7472 14476
rect 7524 14467 7530 14476
rect 7607 14467 7665 14473
rect 7524 14439 7566 14467
rect 7524 14424 7530 14439
rect 7607 14433 7619 14467
rect 7653 14464 7665 14467
rect 7742 14464 7748 14476
rect 7653 14436 7748 14464
rect 7653 14433 7665 14436
rect 7607 14427 7665 14433
rect 7742 14424 7748 14436
rect 7800 14424 7806 14476
rect 9858 14464 9864 14476
rect 9822 14436 9864 14464
rect 9858 14424 9864 14436
rect 9916 14464 9922 14476
rect 10137 14467 10195 14473
rect 10137 14464 10149 14467
rect 9916 14436 10149 14464
rect 9916 14424 9922 14436
rect 10137 14433 10149 14436
rect 10183 14433 10195 14467
rect 10137 14427 10195 14433
rect 10505 14467 10563 14473
rect 10505 14433 10517 14467
rect 10551 14464 10563 14467
rect 11333 14467 11391 14473
rect 10551 14436 10732 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14396 5411 14399
rect 5442 14396 5448 14408
rect 5399 14368 5448 14396
rect 5399 14365 5411 14368
rect 5353 14359 5411 14365
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 6457 14399 6515 14405
rect 6457 14365 6469 14399
rect 6503 14396 6515 14399
rect 7282 14396 7288 14408
rect 6503 14368 7288 14396
rect 6503 14365 6515 14368
rect 6457 14359 6515 14365
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 9122 14396 9128 14408
rect 8352 14368 9128 14396
rect 8352 14356 8358 14368
rect 9122 14356 9128 14368
rect 9180 14396 9186 14408
rect 9401 14399 9459 14405
rect 9401 14396 9413 14399
rect 9180 14368 9413 14396
rect 9180 14356 9186 14368
rect 9401 14365 9413 14368
rect 9447 14396 9459 14399
rect 10597 14399 10655 14405
rect 10597 14396 10609 14399
rect 9447 14368 10609 14396
rect 9447 14365 9459 14368
rect 9401 14359 9459 14365
rect 10597 14365 10609 14368
rect 10643 14365 10655 14399
rect 10597 14359 10655 14365
rect 4246 14220 4252 14272
rect 4304 14260 4310 14272
rect 4709 14263 4767 14269
rect 4709 14260 4721 14263
rect 4304 14232 4721 14260
rect 4304 14220 4310 14232
rect 4709 14229 4721 14232
rect 4755 14229 4767 14263
rect 5460 14260 5488 14356
rect 6638 14288 6644 14340
rect 6696 14328 6702 14340
rect 8110 14328 8116 14340
rect 6696 14300 8116 14328
rect 6696 14288 6702 14300
rect 8110 14288 8116 14300
rect 8168 14288 8174 14340
rect 9490 14288 9496 14340
rect 9548 14328 9554 14340
rect 10704 14328 10732 14436
rect 11333 14433 11345 14467
rect 11379 14464 11391 14467
rect 11698 14464 11704 14476
rect 11379 14436 11704 14464
rect 11379 14433 11391 14436
rect 11333 14427 11391 14433
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 11977 14467 12035 14473
rect 11977 14433 11989 14467
rect 12023 14464 12035 14467
rect 12084 14464 12112 14560
rect 12268 14541 12296 14572
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 12897 14603 12955 14609
rect 12897 14569 12909 14603
rect 12943 14600 12955 14603
rect 13170 14600 13176 14612
rect 12943 14572 13176 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 13906 14560 13912 14612
rect 13964 14560 13970 14612
rect 14182 14560 14188 14612
rect 14240 14560 14246 14612
rect 17402 14560 17408 14612
rect 17460 14600 17466 14612
rect 17681 14603 17739 14609
rect 17681 14600 17693 14603
rect 17460 14572 17693 14600
rect 17460 14560 17466 14572
rect 17681 14569 17693 14572
rect 17727 14569 17739 14603
rect 17681 14563 17739 14569
rect 18414 14560 18420 14612
rect 18472 14560 18478 14612
rect 20162 14560 20168 14612
rect 20220 14560 20226 14612
rect 21085 14603 21143 14609
rect 21085 14569 21097 14603
rect 21131 14569 21143 14603
rect 21085 14563 21143 14569
rect 12161 14535 12219 14541
rect 12161 14501 12173 14535
rect 12207 14532 12219 14535
rect 12253 14535 12311 14541
rect 12253 14532 12265 14535
rect 12207 14504 12265 14532
rect 12207 14501 12219 14504
rect 12161 14495 12219 14501
rect 12253 14501 12265 14504
rect 12299 14501 12311 14535
rect 12253 14495 12311 14501
rect 12526 14492 12532 14544
rect 12584 14495 12590 14544
rect 12989 14535 13047 14541
rect 12989 14501 13001 14535
rect 13035 14532 13047 14535
rect 13078 14532 13084 14544
rect 13035 14504 13084 14532
rect 13035 14501 13047 14504
rect 12989 14495 13047 14501
rect 12584 14492 12596 14495
rect 13078 14492 13084 14504
rect 13136 14492 13142 14544
rect 12538 14489 12596 14492
rect 12023 14436 12112 14464
rect 12023 14433 12035 14436
rect 11977 14427 12035 14433
rect 12434 14424 12440 14476
rect 12492 14424 12498 14476
rect 12538 14455 12550 14489
rect 12584 14455 12596 14489
rect 13924 14473 13952 14560
rect 12538 14449 12596 14455
rect 13173 14467 13231 14473
rect 13173 14433 13185 14467
rect 13219 14464 13231 14467
rect 13909 14467 13967 14473
rect 13219 14436 13308 14464
rect 13219 14433 13231 14436
rect 13173 14427 13231 14433
rect 11422 14356 11428 14408
rect 11480 14356 11486 14408
rect 11606 14356 11612 14408
rect 11664 14396 11670 14408
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 11664 14368 11805 14396
rect 11664 14356 11670 14368
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 12621 14399 12679 14405
rect 12621 14396 12633 14399
rect 11793 14359 11851 14365
rect 11900 14368 12633 14396
rect 9548 14300 10732 14328
rect 9548 14288 9554 14300
rect 10962 14288 10968 14340
rect 11020 14328 11026 14340
rect 11900 14328 11928 14368
rect 12621 14365 12633 14368
rect 12667 14365 12679 14399
rect 12621 14359 12679 14365
rect 13280 14340 13308 14436
rect 13909 14433 13921 14467
rect 13955 14433 13967 14467
rect 13909 14427 13967 14433
rect 14001 14467 14059 14473
rect 14001 14433 14013 14467
rect 14047 14464 14059 14467
rect 14200 14464 14228 14560
rect 16390 14492 16396 14544
rect 16448 14532 16454 14544
rect 19552 14535 19610 14541
rect 16448 14504 18736 14532
rect 16448 14492 16454 14504
rect 18708 14476 18736 14504
rect 19552 14501 19564 14535
rect 19598 14532 19610 14535
rect 20180 14532 20208 14560
rect 19598 14504 20208 14532
rect 21100 14532 21128 14563
rect 21634 14560 21640 14612
rect 21692 14600 21698 14612
rect 22281 14603 22339 14609
rect 22281 14600 22293 14603
rect 21692 14572 22293 14600
rect 21692 14560 21698 14572
rect 22281 14569 22293 14572
rect 22327 14600 22339 14603
rect 22462 14600 22468 14612
rect 22327 14572 22468 14600
rect 22327 14569 22339 14572
rect 22281 14563 22339 14569
rect 22462 14560 22468 14572
rect 22520 14600 22526 14612
rect 22520 14572 22600 14600
rect 22520 14560 22526 14572
rect 21100 14504 21579 14532
rect 19598 14501 19610 14504
rect 19552 14495 19610 14501
rect 14047 14436 14228 14464
rect 17589 14467 17647 14473
rect 14047 14433 14059 14436
rect 14001 14427 14059 14433
rect 17589 14433 17601 14467
rect 17635 14464 17647 14467
rect 17770 14464 17776 14476
rect 17635 14436 17776 14464
rect 17635 14433 17647 14436
rect 17589 14427 17647 14433
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 18690 14424 18696 14476
rect 18748 14464 18754 14476
rect 19702 14464 19708 14476
rect 18748 14436 19708 14464
rect 18748 14424 18754 14436
rect 19702 14424 19708 14436
rect 19760 14464 19766 14476
rect 19797 14467 19855 14473
rect 19797 14464 19809 14467
rect 19760 14436 19809 14464
rect 19760 14424 19766 14436
rect 19797 14433 19809 14436
rect 19843 14433 19855 14467
rect 19797 14427 19855 14433
rect 20809 14467 20867 14473
rect 20809 14433 20821 14467
rect 20855 14433 20867 14467
rect 20809 14427 20867 14433
rect 13633 14399 13691 14405
rect 13633 14365 13645 14399
rect 13679 14396 13691 14399
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13679 14368 13737 14396
rect 13679 14365 13691 14368
rect 13633 14359 13691 14365
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 13725 14359 13783 14365
rect 15838 14356 15844 14408
rect 15896 14396 15902 14408
rect 17865 14399 17923 14405
rect 17865 14396 17877 14399
rect 15896 14368 17877 14396
rect 15896 14356 15902 14368
rect 17865 14365 17877 14368
rect 17911 14396 17923 14399
rect 20824 14396 20852 14427
rect 21450 14424 21456 14476
rect 21508 14424 21514 14476
rect 21551 14464 21579 14504
rect 21744 14504 22416 14532
rect 21744 14464 21772 14504
rect 21551 14436 21772 14464
rect 21913 14467 21971 14473
rect 21913 14462 21925 14467
rect 21836 14434 21925 14462
rect 20990 14396 20996 14408
rect 17911 14368 18000 14396
rect 20824 14368 20996 14396
rect 17911 14365 17923 14368
rect 17865 14359 17923 14365
rect 11020 14300 11928 14328
rect 12253 14331 12311 14337
rect 11020 14288 11026 14300
rect 12253 14297 12265 14331
rect 12299 14328 12311 14331
rect 13262 14328 13268 14340
rect 12299 14300 13268 14328
rect 12299 14297 12311 14300
rect 12253 14291 12311 14297
rect 13262 14288 13268 14300
rect 13320 14288 13326 14340
rect 7190 14260 7196 14272
rect 5460 14232 7196 14260
rect 4709 14223 4767 14229
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 7834 14220 7840 14272
rect 7892 14220 7898 14272
rect 7926 14220 7932 14272
rect 7984 14220 7990 14272
rect 10042 14220 10048 14272
rect 10100 14220 10106 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 12713 14263 12771 14269
rect 12713 14260 12725 14263
rect 11940 14232 12725 14260
rect 11940 14220 11946 14232
rect 12713 14229 12725 14232
rect 12759 14229 12771 14263
rect 12713 14223 12771 14229
rect 12805 14263 12863 14269
rect 12805 14229 12817 14263
rect 12851 14260 12863 14263
rect 13449 14263 13507 14269
rect 13449 14260 13461 14263
rect 12851 14232 13461 14260
rect 12851 14229 12863 14232
rect 12805 14223 12863 14229
rect 13449 14229 13461 14232
rect 13495 14260 13507 14263
rect 13722 14260 13728 14272
rect 13495 14232 13728 14260
rect 13495 14229 13507 14232
rect 13449 14223 13507 14229
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 13814 14220 13820 14272
rect 13872 14220 13878 14272
rect 16758 14220 16764 14272
rect 16816 14260 16822 14272
rect 17221 14263 17279 14269
rect 17221 14260 17233 14263
rect 16816 14232 17233 14260
rect 16816 14220 16822 14232
rect 17221 14229 17233 14232
rect 17267 14229 17279 14263
rect 17972 14260 18000 14368
rect 20990 14356 20996 14368
rect 21048 14356 21054 14408
rect 21088 14399 21146 14405
rect 21088 14365 21100 14399
rect 21134 14396 21146 14399
rect 21134 14368 21496 14396
rect 21134 14365 21146 14368
rect 21088 14359 21146 14365
rect 21468 14340 21496 14368
rect 21542 14356 21548 14408
rect 21600 14356 21606 14408
rect 21836 14396 21864 14434
rect 21913 14433 21925 14434
rect 21959 14433 21971 14467
rect 21913 14427 21971 14433
rect 22094 14424 22100 14476
rect 22152 14424 22158 14476
rect 22388 14473 22416 14504
rect 22572 14473 22600 14572
rect 22373 14467 22431 14473
rect 22373 14433 22385 14467
rect 22419 14433 22431 14467
rect 22373 14427 22431 14433
rect 22557 14467 22615 14473
rect 22557 14433 22569 14467
rect 22603 14433 22615 14467
rect 22557 14427 22615 14433
rect 21652 14368 21864 14396
rect 21450 14288 21456 14340
rect 21508 14288 21514 14340
rect 19426 14260 19432 14272
rect 17972 14232 19432 14260
rect 17221 14223 17279 14229
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 20901 14263 20959 14269
rect 20901 14229 20913 14263
rect 20947 14260 20959 14263
rect 21174 14260 21180 14272
rect 20947 14232 21180 14260
rect 20947 14229 20959 14232
rect 20901 14223 20959 14229
rect 21174 14220 21180 14232
rect 21232 14260 21238 14272
rect 21652 14260 21680 14368
rect 21836 14300 22692 14328
rect 21836 14269 21864 14300
rect 22664 14272 22692 14300
rect 21232 14232 21680 14260
rect 21821 14263 21879 14269
rect 21232 14220 21238 14232
rect 21821 14229 21833 14263
rect 21867 14229 21879 14263
rect 21821 14223 21879 14229
rect 22097 14263 22155 14269
rect 22097 14229 22109 14263
rect 22143 14260 22155 14263
rect 22186 14260 22192 14272
rect 22143 14232 22192 14260
rect 22143 14229 22155 14232
rect 22097 14223 22155 14229
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 22462 14220 22468 14272
rect 22520 14220 22526 14272
rect 22646 14220 22652 14272
rect 22704 14220 22710 14272
rect 552 14170 23368 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 23368 14170
rect 552 14096 23368 14118
rect 5718 14016 5724 14068
rect 5776 14016 5782 14068
rect 7190 14016 7196 14068
rect 7248 14016 7254 14068
rect 9585 14059 9643 14065
rect 9585 14025 9597 14059
rect 9631 14056 9643 14059
rect 9858 14056 9864 14068
rect 9631 14028 9864 14056
rect 9631 14025 9643 14028
rect 9585 14019 9643 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 11422 14016 11428 14068
rect 11480 14056 11486 14068
rect 11609 14059 11667 14065
rect 11609 14056 11621 14059
rect 11480 14028 11621 14056
rect 11480 14016 11486 14028
rect 11609 14025 11621 14028
rect 11655 14025 11667 14059
rect 12434 14056 12440 14068
rect 11609 14019 11667 14025
rect 12406 14016 12440 14056
rect 12492 14016 12498 14068
rect 13814 14016 13820 14068
rect 13872 14016 13878 14068
rect 16758 14056 16764 14068
rect 16592 14028 16764 14056
rect 7208 13988 7236 14016
rect 10226 13988 10232 14000
rect 7208 13960 10232 13988
rect 10226 13948 10232 13960
rect 10284 13948 10290 14000
rect 7653 13923 7711 13929
rect 7653 13889 7665 13923
rect 7699 13920 7711 13923
rect 7926 13920 7932 13932
rect 7699 13892 7932 13920
rect 7699 13889 7711 13892
rect 7653 13883 7711 13889
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 8202 13880 8208 13932
rect 8260 13920 8266 13932
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 8260 13892 8493 13920
rect 8260 13880 8266 13892
rect 8481 13889 8493 13892
rect 8527 13920 8539 13923
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 8527 13892 9505 13920
rect 8527 13889 8539 13892
rect 8481 13883 8539 13889
rect 9493 13889 9505 13892
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 11422 13880 11428 13932
rect 11480 13920 11486 13932
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11480 13892 11805 13920
rect 11480 13880 11486 13892
rect 11793 13889 11805 13892
rect 11839 13920 11851 13923
rect 12406 13920 12434 14016
rect 11839 13892 12434 13920
rect 11839 13889 11851 13892
rect 11793 13883 11851 13889
rect 13262 13880 13268 13932
rect 13320 13920 13326 13932
rect 13633 13923 13691 13929
rect 13633 13920 13645 13923
rect 13320 13892 13645 13920
rect 13320 13880 13326 13892
rect 13633 13889 13645 13892
rect 13679 13889 13691 13923
rect 13832 13920 13860 14016
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 13832 13892 14289 13920
rect 13633 13883 13691 13889
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 15194 13880 15200 13932
rect 15252 13920 15258 13932
rect 15657 13923 15715 13929
rect 15657 13920 15669 13923
rect 15252 13892 15669 13920
rect 15252 13880 15258 13892
rect 15657 13889 15669 13892
rect 15703 13889 15715 13923
rect 15657 13883 15715 13889
rect 15838 13880 15844 13932
rect 15896 13880 15902 13932
rect 16390 13880 16396 13932
rect 16448 13880 16454 13932
rect 4341 13855 4399 13861
rect 4341 13821 4353 13855
rect 4387 13852 4399 13855
rect 4430 13852 4436 13864
rect 4387 13824 4436 13852
rect 4387 13821 4399 13824
rect 4341 13815 4399 13821
rect 4430 13812 4436 13824
rect 4488 13812 4494 13864
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 7561 13855 7619 13861
rect 7561 13852 7573 13855
rect 6788 13824 7573 13852
rect 6788 13812 6794 13824
rect 7561 13821 7573 13824
rect 7607 13821 7619 13855
rect 7561 13815 7619 13821
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 8352 13824 8401 13852
rect 8352 13812 8358 13824
rect 8389 13821 8401 13824
rect 8435 13821 8447 13855
rect 8389 13815 8447 13821
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 4154 13744 4160 13796
rect 4212 13784 4218 13796
rect 4586 13787 4644 13793
rect 4586 13784 4598 13787
rect 4212 13756 4598 13784
rect 4212 13744 4218 13756
rect 4586 13753 4598 13756
rect 4632 13753 4644 13787
rect 4586 13747 4644 13753
rect 8588 13728 8616 13815
rect 9398 13812 9404 13864
rect 9456 13812 9462 13864
rect 11241 13855 11299 13861
rect 11241 13852 11253 13855
rect 10060 13824 11253 13852
rect 10060 13796 10088 13824
rect 11241 13821 11253 13824
rect 11287 13821 11299 13855
rect 11241 13815 11299 13821
rect 11517 13855 11575 13861
rect 11517 13821 11529 13855
rect 11563 13852 11575 13855
rect 11698 13852 11704 13864
rect 11563 13824 11704 13852
rect 11563 13821 11575 13824
rect 11517 13815 11575 13821
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 13078 13812 13084 13864
rect 13136 13852 13142 13864
rect 13136 13824 13676 13852
rect 13136 13812 13142 13824
rect 10042 13744 10048 13796
rect 10100 13744 10106 13796
rect 10962 13744 10968 13796
rect 11020 13784 11026 13796
rect 11057 13787 11115 13793
rect 11057 13784 11069 13787
rect 11020 13756 11069 13784
rect 11020 13744 11026 13756
rect 11057 13753 11069 13756
rect 11103 13753 11115 13787
rect 13648 13784 13676 13824
rect 13722 13812 13728 13864
rect 13780 13812 13786 13864
rect 14369 13855 14427 13861
rect 14369 13852 14381 13855
rect 13832 13824 14381 13852
rect 13832 13784 13860 13824
rect 14369 13821 14381 13824
rect 14415 13821 14427 13855
rect 14369 13815 14427 13821
rect 16022 13812 16028 13864
rect 16080 13812 16086 13864
rect 13648 13756 13860 13784
rect 11057 13747 11115 13753
rect 16114 13744 16120 13796
rect 16172 13784 16178 13796
rect 16408 13784 16436 13880
rect 16485 13855 16543 13861
rect 16485 13821 16497 13855
rect 16531 13852 16543 13855
rect 16592 13852 16620 14028
rect 16758 14016 16764 14028
rect 16816 14016 16822 14068
rect 17034 14016 17040 14068
rect 17092 14056 17098 14068
rect 17092 14028 17724 14056
rect 17092 14016 17098 14028
rect 16669 13991 16727 13997
rect 16669 13957 16681 13991
rect 16715 13957 16727 13991
rect 17696 13988 17724 14028
rect 17770 14016 17776 14068
rect 17828 14056 17834 14068
rect 18141 14059 18199 14065
rect 18141 14056 18153 14059
rect 17828 14028 18153 14056
rect 17828 14016 17834 14028
rect 18141 14025 18153 14028
rect 18187 14025 18199 14059
rect 18141 14019 18199 14025
rect 19426 14016 19432 14068
rect 19484 14056 19490 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19484 14028 19533 14056
rect 19484 14016 19490 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 21450 14016 21456 14068
rect 21508 14056 21514 14068
rect 22186 14056 22192 14068
rect 21508 14028 22192 14056
rect 21508 14016 21514 14028
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 19153 13991 19211 13997
rect 19153 13988 19165 13991
rect 17696 13960 19165 13988
rect 16669 13951 16727 13957
rect 19153 13957 19165 13960
rect 19199 13988 19211 13991
rect 20714 13988 20720 14000
rect 19199 13960 20720 13988
rect 19199 13957 19211 13960
rect 19153 13951 19211 13957
rect 16684 13920 16712 13951
rect 20714 13948 20720 13960
rect 20772 13948 20778 14000
rect 20809 13923 20867 13929
rect 16684 13892 16896 13920
rect 16761 13855 16819 13861
rect 16761 13852 16773 13855
rect 16531 13824 16620 13852
rect 16684 13824 16773 13852
rect 16531 13821 16543 13824
rect 16485 13815 16543 13821
rect 16684 13784 16712 13824
rect 16761 13821 16773 13824
rect 16807 13821 16819 13855
rect 16868 13852 16896 13892
rect 20809 13889 20821 13923
rect 20855 13920 20867 13923
rect 21174 13920 21180 13932
rect 20855 13892 21180 13920
rect 20855 13889 20867 13892
rect 20809 13883 20867 13889
rect 21174 13880 21180 13892
rect 21232 13880 21238 13932
rect 21450 13880 21456 13932
rect 21508 13880 21514 13932
rect 17017 13855 17075 13861
rect 17017 13852 17029 13855
rect 16868 13824 17029 13852
rect 16761 13815 16819 13821
rect 17017 13821 17029 13824
rect 17063 13821 17075 13855
rect 17017 13815 17075 13821
rect 18969 13855 19027 13861
rect 18969 13821 18981 13855
rect 19015 13852 19027 13855
rect 19334 13852 19340 13864
rect 19015 13824 19340 13852
rect 19015 13821 19027 13824
rect 18969 13815 19027 13821
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 19429 13855 19487 13861
rect 19429 13821 19441 13855
rect 19475 13852 19487 13855
rect 19518 13852 19524 13864
rect 19475 13824 19524 13852
rect 19475 13821 19487 13824
rect 19429 13815 19487 13821
rect 19518 13812 19524 13824
rect 19576 13852 19582 13864
rect 20346 13852 20352 13864
rect 19576 13824 20352 13852
rect 19576 13812 19582 13824
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 20530 13812 20536 13864
rect 20588 13852 20594 13864
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20588 13824 20637 13852
rect 20588 13812 20594 13824
rect 20625 13821 20637 13824
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 20990 13812 20996 13864
rect 21048 13852 21054 13864
rect 21085 13855 21143 13861
rect 21085 13852 21097 13855
rect 21048 13824 21097 13852
rect 21048 13812 21054 13824
rect 21085 13821 21097 13824
rect 21131 13852 21143 13855
rect 22094 13852 22100 13864
rect 21131 13824 22100 13852
rect 21131 13821 21143 13824
rect 21085 13815 21143 13821
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 16172 13756 16712 13784
rect 16172 13744 16178 13756
rect 20438 13744 20444 13796
rect 20496 13744 20502 13796
rect 7929 13719 7987 13725
rect 7929 13685 7941 13719
rect 7975 13716 7987 13719
rect 8570 13716 8576 13728
rect 7975 13688 8576 13716
rect 7975 13685 7987 13688
rect 7929 13679 7987 13685
rect 8570 13676 8576 13688
rect 8628 13676 8634 13728
rect 9766 13676 9772 13728
rect 9824 13676 9830 13728
rect 11790 13676 11796 13728
rect 11848 13676 11854 13728
rect 14090 13676 14096 13728
rect 14148 13676 14154 13728
rect 14737 13719 14795 13725
rect 14737 13685 14749 13719
rect 14783 13716 14795 13719
rect 14826 13716 14832 13728
rect 14783 13688 14832 13716
rect 14783 13685 14795 13688
rect 14737 13679 14795 13685
rect 14826 13676 14832 13688
rect 14884 13676 14890 13728
rect 15194 13676 15200 13728
rect 15252 13676 15258 13728
rect 15565 13719 15623 13725
rect 15565 13685 15577 13719
rect 15611 13716 15623 13719
rect 15930 13716 15936 13728
rect 15611 13688 15936 13716
rect 15611 13685 15623 13688
rect 15565 13679 15623 13685
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 16206 13676 16212 13728
rect 16264 13676 16270 13728
rect 552 13626 23368 13648
rect 552 13574 19022 13626
rect 19074 13574 19086 13626
rect 19138 13574 19150 13626
rect 19202 13574 19214 13626
rect 19266 13574 19278 13626
rect 19330 13574 23368 13626
rect 552 13552 23368 13574
rect 3881 13515 3939 13521
rect 3881 13481 3893 13515
rect 3927 13512 3939 13515
rect 4062 13512 4068 13524
rect 3927 13484 4068 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4157 13515 4215 13521
rect 4157 13481 4169 13515
rect 4203 13481 4215 13515
rect 4157 13475 4215 13481
rect 4172 13444 4200 13475
rect 5626 13472 5632 13524
rect 5684 13512 5690 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 5684 13484 6285 13512
rect 5684 13472 5690 13484
rect 6273 13481 6285 13484
rect 6319 13481 6331 13515
rect 6273 13475 6331 13481
rect 8570 13472 8576 13524
rect 8628 13472 8634 13524
rect 17034 13512 17040 13524
rect 12406 13484 17040 13512
rect 4494 13447 4552 13453
rect 4494 13444 4506 13447
rect 4172 13416 4506 13444
rect 4494 13413 4506 13416
rect 4540 13413 4552 13447
rect 4494 13407 4552 13413
rect 5350 13404 5356 13456
rect 5408 13444 5414 13456
rect 6181 13447 6239 13453
rect 6181 13444 6193 13447
rect 5408 13416 6193 13444
rect 5408 13404 5414 13416
rect 6181 13413 6193 13416
rect 6227 13413 6239 13447
rect 6181 13407 6239 13413
rect 3697 13379 3755 13385
rect 3697 13345 3709 13379
rect 3743 13345 3755 13379
rect 3697 13339 3755 13345
rect 3973 13379 4031 13385
rect 3973 13345 3985 13379
rect 4019 13376 4031 13379
rect 6822 13376 6828 13388
rect 4019 13348 5856 13376
rect 4019 13345 4031 13348
rect 3973 13339 4031 13345
rect 3712 13308 3740 13339
rect 4154 13308 4160 13320
rect 3712 13280 4160 13308
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13277 4307 13311
rect 4249 13271 4307 13277
rect 4264 13172 4292 13271
rect 5828 13249 5856 13348
rect 6472 13348 6828 13376
rect 6472 13317 6500 13348
rect 6822 13336 6828 13348
rect 6880 13376 6886 13388
rect 7926 13376 7932 13388
rect 6880 13348 7932 13376
rect 6880 13336 6886 13348
rect 7926 13336 7932 13348
rect 7984 13336 7990 13388
rect 8202 13336 8208 13388
rect 8260 13336 8266 13388
rect 8386 13336 8392 13388
rect 8444 13336 8450 13388
rect 8588 13376 8616 13472
rect 12406 13444 12434 13484
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 19521 13515 19579 13521
rect 19521 13481 19533 13515
rect 19567 13512 19579 13515
rect 19567 13484 20208 13512
rect 19567 13481 19579 13484
rect 19521 13475 19579 13481
rect 10244 13416 12434 13444
rect 14568 13416 16160 13444
rect 10244 13388 10272 13416
rect 8665 13379 8723 13385
rect 8665 13376 8677 13379
rect 8588 13348 8677 13376
rect 8665 13345 8677 13348
rect 8711 13345 8723 13379
rect 8665 13339 8723 13345
rect 8757 13379 8815 13385
rect 8757 13345 8769 13379
rect 8803 13345 8815 13379
rect 8757 13339 8815 13345
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 8294 13308 8300 13320
rect 7432 13280 8300 13308
rect 7432 13268 7438 13280
rect 8294 13268 8300 13280
rect 8352 13308 8358 13320
rect 8772 13308 8800 13339
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 9824 13348 10149 13376
rect 9824 13336 9830 13348
rect 10137 13345 10149 13348
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 10226 13336 10232 13388
rect 10284 13336 10290 13388
rect 10597 13379 10655 13385
rect 10597 13345 10609 13379
rect 10643 13345 10655 13379
rect 10597 13339 10655 13345
rect 10781 13379 10839 13385
rect 10781 13345 10793 13379
rect 10827 13376 10839 13379
rect 10962 13376 10968 13388
rect 10827 13348 10968 13376
rect 10827 13345 10839 13348
rect 10781 13339 10839 13345
rect 8352 13280 8800 13308
rect 8352 13268 8358 13280
rect 10042 13268 10048 13320
rect 10100 13268 10106 13320
rect 10318 13268 10324 13320
rect 10376 13268 10382 13320
rect 5813 13243 5871 13249
rect 5813 13209 5825 13243
rect 5859 13209 5871 13243
rect 5813 13203 5871 13209
rect 8067 13243 8125 13249
rect 8067 13209 8079 13243
rect 8113 13240 8125 13243
rect 8481 13243 8539 13249
rect 8481 13240 8493 13243
rect 8113 13212 8493 13240
rect 8113 13209 8125 13212
rect 8067 13203 8125 13209
rect 8481 13209 8493 13212
rect 8527 13209 8539 13243
rect 10060 13240 10088 13268
rect 10612 13240 10640 13339
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 11164 13385 11192 13416
rect 14568 13388 14596 13416
rect 16132 13388 16160 13416
rect 16206 13404 16212 13456
rect 16264 13444 16270 13456
rect 16362 13447 16420 13453
rect 16362 13444 16374 13447
rect 16264 13416 16374 13444
rect 16264 13404 16270 13416
rect 16362 13413 16374 13416
rect 16408 13413 16420 13447
rect 16362 13407 16420 13413
rect 19794 13404 19800 13456
rect 19852 13404 19858 13456
rect 19889 13447 19947 13453
rect 19889 13413 19901 13447
rect 19935 13444 19947 13447
rect 19935 13416 20024 13444
rect 19935 13413 19947 13416
rect 19889 13407 19947 13413
rect 11149 13379 11207 13385
rect 11149 13345 11161 13379
rect 11195 13345 11207 13379
rect 11149 13339 11207 13345
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13376 11299 13379
rect 11422 13376 11428 13388
rect 11287 13348 11428 13376
rect 11287 13345 11299 13348
rect 11241 13339 11299 13345
rect 11422 13336 11428 13348
rect 11480 13336 11486 13388
rect 11974 13336 11980 13388
rect 12032 13336 12038 13388
rect 14550 13336 14556 13388
rect 14608 13336 14614 13388
rect 14820 13379 14878 13385
rect 14820 13345 14832 13379
rect 14866 13376 14878 13379
rect 15102 13376 15108 13388
rect 14866 13348 15108 13376
rect 14866 13345 14878 13348
rect 14820 13339 14878 13345
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 16114 13336 16120 13388
rect 16172 13336 16178 13388
rect 19153 13379 19211 13385
rect 19153 13376 19165 13379
rect 18800 13348 19165 13376
rect 11054 13268 11060 13320
rect 11112 13268 11118 13320
rect 11333 13311 11391 13317
rect 11333 13277 11345 13311
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 10060 13212 10640 13240
rect 10689 13243 10747 13249
rect 8481 13203 8539 13209
rect 10689 13209 10701 13243
rect 10735 13240 10747 13243
rect 11348 13240 11376 13271
rect 11790 13268 11796 13320
rect 11848 13308 11854 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11848 13280 11897 13308
rect 11848 13268 11854 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 18800 13252 18828 13348
rect 19153 13345 19165 13348
rect 19199 13345 19211 13379
rect 19153 13339 19211 13345
rect 19168 13308 19196 13339
rect 19334 13336 19340 13388
rect 19392 13376 19398 13388
rect 19613 13379 19671 13385
rect 19613 13376 19625 13379
rect 19392 13348 19625 13376
rect 19392 13336 19398 13348
rect 19613 13345 19625 13348
rect 19659 13376 19671 13379
rect 19812 13376 19840 13404
rect 19996 13385 20024 13416
rect 20180 13385 20208 13484
rect 20530 13472 20536 13524
rect 20588 13472 20594 13524
rect 20714 13472 20720 13524
rect 20772 13512 20778 13524
rect 21427 13515 21485 13521
rect 21427 13512 21439 13515
rect 20772 13484 21439 13512
rect 20772 13472 20778 13484
rect 21427 13481 21439 13484
rect 21473 13481 21485 13515
rect 21427 13475 21485 13481
rect 20548 13444 20576 13472
rect 20548 13416 20760 13444
rect 19659 13348 19840 13376
rect 19981 13379 20039 13385
rect 19659 13345 19671 13348
rect 19613 13339 19671 13345
rect 19981 13345 19993 13379
rect 20027 13345 20039 13379
rect 19981 13339 20039 13345
rect 20165 13379 20223 13385
rect 20165 13345 20177 13379
rect 20211 13376 20223 13379
rect 20438 13376 20444 13388
rect 20211 13348 20444 13376
rect 20211 13345 20223 13348
rect 20165 13339 20223 13345
rect 20438 13336 20444 13348
rect 20496 13376 20502 13388
rect 20732 13385 20760 13416
rect 21174 13404 21180 13456
rect 21232 13444 21238 13456
rect 21637 13447 21695 13453
rect 21637 13444 21649 13447
rect 21232 13416 21649 13444
rect 21232 13404 21238 13416
rect 21637 13413 21649 13416
rect 21683 13413 21695 13447
rect 21637 13407 21695 13413
rect 20533 13379 20591 13385
rect 20533 13376 20545 13379
rect 20496 13348 20545 13376
rect 20496 13336 20502 13348
rect 20533 13345 20545 13348
rect 20579 13345 20591 13379
rect 20533 13339 20591 13345
rect 20717 13379 20775 13385
rect 20717 13345 20729 13379
rect 20763 13345 20775 13379
rect 20717 13339 20775 13345
rect 21266 13336 21272 13388
rect 21324 13336 21330 13388
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19168 13280 19717 13308
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13277 19947 13311
rect 19889 13271 19947 13277
rect 10735 13212 11376 13240
rect 12345 13243 12403 13249
rect 10735 13209 10747 13212
rect 10689 13203 10747 13209
rect 12345 13209 12357 13243
rect 12391 13240 12403 13243
rect 12894 13240 12900 13252
rect 12391 13212 12900 13240
rect 12391 13209 12403 13212
rect 12345 13203 12403 13209
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 18782 13200 18788 13252
rect 18840 13200 18846 13252
rect 19904 13240 19932 13271
rect 19168 13212 19932 13240
rect 4522 13172 4528 13184
rect 4264 13144 4528 13172
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 8294 13132 8300 13184
rect 8352 13132 8358 13184
rect 9858 13132 9864 13184
rect 9916 13132 9922 13184
rect 11514 13132 11520 13184
rect 11572 13132 11578 13184
rect 15930 13132 15936 13184
rect 15988 13132 15994 13184
rect 17497 13175 17555 13181
rect 17497 13141 17509 13175
rect 17543 13172 17555 13175
rect 17586 13172 17592 13184
rect 17543 13144 17592 13172
rect 17543 13141 17555 13144
rect 17497 13135 17555 13141
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 18414 13132 18420 13184
rect 18472 13172 18478 13184
rect 19168 13181 19196 13212
rect 20806 13200 20812 13252
rect 20864 13240 20870 13252
rect 21284 13240 21312 13336
rect 20864 13212 21496 13240
rect 20864 13200 20870 13212
rect 19153 13175 19211 13181
rect 19153 13172 19165 13175
rect 18472 13144 19165 13172
rect 18472 13132 18478 13144
rect 19153 13141 19165 13144
rect 19199 13141 19211 13175
rect 19153 13135 19211 13141
rect 20070 13132 20076 13184
rect 20128 13132 20134 13184
rect 21266 13132 21272 13184
rect 21324 13132 21330 13184
rect 21468 13181 21496 13212
rect 21453 13175 21511 13181
rect 21453 13141 21465 13175
rect 21499 13141 21511 13175
rect 21453 13135 21511 13141
rect 552 13082 23368 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 23368 13082
rect 552 13008 23368 13030
rect 8294 12928 8300 12980
rect 8352 12928 8358 12980
rect 10318 12928 10324 12980
rect 10376 12968 10382 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10376 12940 10425 12968
rect 10376 12928 10382 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 15102 12928 15108 12980
rect 15160 12968 15166 12980
rect 15197 12971 15255 12977
rect 15197 12968 15209 12971
rect 15160 12940 15209 12968
rect 15160 12928 15166 12940
rect 15197 12937 15209 12940
rect 15243 12937 15255 12971
rect 15197 12931 15255 12937
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 16393 12971 16451 12977
rect 16393 12968 16405 12971
rect 16080 12940 16405 12968
rect 16080 12928 16086 12940
rect 16393 12937 16405 12940
rect 16439 12937 16451 12971
rect 16393 12931 16451 12937
rect 17589 12971 17647 12977
rect 17589 12937 17601 12971
rect 17635 12968 17647 12971
rect 17678 12968 17684 12980
rect 17635 12940 17684 12968
rect 17635 12937 17647 12940
rect 17589 12931 17647 12937
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 20714 12928 20720 12980
rect 20772 12928 20778 12980
rect 21450 12928 21456 12980
rect 21508 12928 21514 12980
rect 4246 12724 4252 12776
rect 4304 12724 4310 12776
rect 4522 12724 4528 12776
rect 4580 12764 4586 12776
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 4580 12736 6837 12764
rect 4580 12724 4586 12736
rect 6825 12733 6837 12736
rect 6871 12764 6883 12767
rect 8312 12764 8340 12928
rect 14277 12903 14335 12909
rect 14277 12869 14289 12903
rect 14323 12900 14335 12903
rect 15286 12900 15292 12912
rect 14323 12872 15292 12900
rect 14323 12869 14335 12872
rect 14277 12863 14335 12869
rect 15286 12860 15292 12872
rect 15344 12860 15350 12912
rect 17773 12903 17831 12909
rect 15396 12872 15884 12900
rect 13725 12835 13783 12841
rect 13725 12801 13737 12835
rect 13771 12801 13783 12835
rect 13725 12795 13783 12801
rect 13817 12835 13875 12841
rect 13817 12801 13829 12835
rect 13863 12832 13875 12835
rect 14090 12832 14096 12844
rect 13863 12804 14096 12832
rect 13863 12801 13875 12804
rect 13817 12795 13875 12801
rect 9502 12767 9560 12773
rect 9502 12764 9514 12767
rect 6871 12736 7604 12764
rect 8312 12736 9514 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 4770 12699 4828 12705
rect 4770 12696 4782 12699
rect 4448 12668 4782 12696
rect 4448 12637 4476 12668
rect 4770 12665 4782 12668
rect 4816 12665 4828 12699
rect 4770 12659 4828 12665
rect 7092 12699 7150 12705
rect 7092 12665 7104 12699
rect 7138 12696 7150 12699
rect 7466 12696 7472 12708
rect 7138 12668 7472 12696
rect 7138 12665 7150 12668
rect 7092 12659 7150 12665
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 7576 12696 7604 12736
rect 9502 12733 9514 12736
rect 9548 12733 9560 12767
rect 9502 12727 9560 12733
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12733 9827 12767
rect 9769 12727 9827 12733
rect 10597 12767 10655 12773
rect 10597 12733 10609 12767
rect 10643 12733 10655 12767
rect 10597 12727 10655 12733
rect 9398 12696 9404 12708
rect 7576 12668 9404 12696
rect 9398 12656 9404 12668
rect 9456 12696 9462 12708
rect 9784 12696 9812 12727
rect 9456 12668 9812 12696
rect 9456 12656 9462 12668
rect 9950 12656 9956 12708
rect 10008 12696 10014 12708
rect 10612 12696 10640 12727
rect 10778 12724 10784 12776
rect 10836 12724 10842 12776
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12764 11759 12767
rect 13740 12764 13768 12795
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 15013 12835 15071 12841
rect 15013 12832 15025 12835
rect 14660 12804 15025 12832
rect 13906 12764 13912 12776
rect 11747 12736 12434 12764
rect 13740 12736 13912 12764
rect 11747 12733 11759 12736
rect 11701 12727 11759 12733
rect 11330 12696 11336 12708
rect 10008 12668 11336 12696
rect 10008 12656 10014 12668
rect 11330 12656 11336 12668
rect 11388 12696 11394 12708
rect 12406 12696 12434 12736
rect 13906 12724 13912 12736
rect 13964 12764 13970 12776
rect 14660 12764 14688 12804
rect 15013 12801 15025 12804
rect 15059 12832 15071 12835
rect 15396 12832 15424 12872
rect 15856 12844 15884 12872
rect 17773 12869 17785 12903
rect 17819 12900 17831 12903
rect 17819 12872 18828 12900
rect 17819 12869 17831 12872
rect 17773 12863 17831 12869
rect 18800 12844 18828 12872
rect 15059 12804 15424 12832
rect 15059 12801 15071 12804
rect 15013 12795 15071 12801
rect 15470 12792 15476 12844
rect 15528 12792 15534 12844
rect 15838 12792 15844 12844
rect 15896 12792 15902 12844
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12832 17555 12835
rect 17543 12804 17816 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 13964 12736 14688 12764
rect 14737 12767 14795 12773
rect 13964 12724 13970 12736
rect 14737 12733 14749 12767
rect 14783 12764 14795 12767
rect 15102 12764 15108 12776
rect 14783 12736 15108 12764
rect 14783 12733 14795 12736
rect 14737 12727 14795 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15381 12767 15439 12773
rect 15381 12764 15393 12767
rect 15252 12736 15393 12764
rect 15252 12724 15258 12736
rect 15381 12733 15393 12736
rect 15427 12733 15439 12767
rect 15488 12764 15516 12792
rect 17788 12776 17816 12804
rect 18782 12792 18788 12844
rect 18840 12792 18846 12844
rect 19245 12835 19303 12841
rect 19245 12801 19257 12835
rect 19291 12832 19303 12835
rect 19426 12832 19432 12844
rect 19291 12804 19432 12832
rect 19291 12801 19303 12804
rect 19245 12795 19303 12801
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 15933 12767 15991 12773
rect 15933 12764 15945 12767
rect 15488 12736 15945 12764
rect 15381 12727 15439 12733
rect 15933 12733 15945 12736
rect 15979 12733 15991 12767
rect 15933 12727 15991 12733
rect 16025 12767 16083 12773
rect 16025 12733 16037 12767
rect 16071 12764 16083 12767
rect 16942 12764 16948 12776
rect 16071 12736 16948 12764
rect 16071 12733 16083 12736
rect 16025 12727 16083 12733
rect 16942 12724 16948 12736
rect 17000 12764 17006 12776
rect 17586 12764 17592 12776
rect 17000 12736 17592 12764
rect 17000 12724 17006 12736
rect 17586 12724 17592 12736
rect 17644 12724 17650 12776
rect 17770 12724 17776 12776
rect 17828 12724 17834 12776
rect 18877 12767 18935 12773
rect 18877 12733 18889 12767
rect 18923 12764 18935 12767
rect 19334 12764 19340 12776
rect 18923 12736 19340 12764
rect 18923 12733 18935 12736
rect 18877 12727 18935 12733
rect 19334 12724 19340 12736
rect 19392 12724 19398 12776
rect 20732 12773 20760 12928
rect 20990 12860 20996 12912
rect 21048 12860 21054 12912
rect 21361 12835 21419 12841
rect 21361 12801 21373 12835
rect 21407 12832 21419 12835
rect 21468 12832 21496 12928
rect 21729 12903 21787 12909
rect 21729 12869 21741 12903
rect 21775 12900 21787 12903
rect 22094 12900 22100 12912
rect 21775 12872 22100 12900
rect 21775 12869 21787 12872
rect 21729 12863 21787 12869
rect 22094 12860 22100 12872
rect 22152 12860 22158 12912
rect 21407 12804 21496 12832
rect 22189 12835 22247 12841
rect 21407 12801 21419 12804
rect 21361 12795 21419 12801
rect 22189 12801 22201 12835
rect 22235 12832 22247 12835
rect 22462 12832 22468 12844
rect 22235 12804 22468 12832
rect 22235 12801 22247 12804
rect 22189 12795 22247 12801
rect 22462 12792 22468 12804
rect 22520 12792 22526 12844
rect 22646 12792 22652 12844
rect 22704 12792 22710 12844
rect 20717 12767 20775 12773
rect 20717 12733 20729 12767
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 20806 12724 20812 12776
rect 20864 12724 20870 12776
rect 20993 12767 21051 12773
rect 20993 12733 21005 12767
rect 21039 12764 21051 12767
rect 21174 12764 21180 12776
rect 21039 12736 21180 12764
rect 21039 12733 21051 12736
rect 20993 12727 21051 12733
rect 21174 12724 21180 12736
rect 21232 12724 21238 12776
rect 21450 12724 21456 12776
rect 21508 12724 21514 12776
rect 21726 12724 21732 12776
rect 21784 12764 21790 12776
rect 22097 12767 22155 12773
rect 22097 12764 22109 12767
rect 21784 12736 22109 12764
rect 21784 12724 21790 12736
rect 22097 12733 22109 12736
rect 22143 12733 22155 12767
rect 22097 12727 22155 12733
rect 22738 12724 22744 12776
rect 22796 12724 22802 12776
rect 11388 12668 11560 12696
rect 12406 12668 14504 12696
rect 11388 12656 11394 12668
rect 4433 12631 4491 12637
rect 4433 12597 4445 12631
rect 4479 12597 4491 12631
rect 4433 12591 4491 12597
rect 5902 12588 5908 12640
rect 5960 12588 5966 12640
rect 8202 12588 8208 12640
rect 8260 12588 8266 12640
rect 8389 12631 8447 12637
rect 8389 12597 8401 12631
rect 8435 12628 8447 12631
rect 8478 12628 8484 12640
rect 8435 12600 8484 12628
rect 8435 12597 8447 12600
rect 8389 12591 8447 12597
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 11532 12637 11560 12668
rect 11517 12631 11575 12637
rect 11517 12597 11529 12631
rect 11563 12597 11575 12631
rect 11517 12591 11575 12597
rect 13906 12588 13912 12640
rect 13964 12588 13970 12640
rect 14366 12588 14372 12640
rect 14424 12588 14430 12640
rect 14476 12628 14504 12668
rect 14826 12656 14832 12708
rect 14884 12656 14890 12708
rect 17218 12656 17224 12708
rect 17276 12696 17282 12708
rect 17313 12699 17371 12705
rect 17313 12696 17325 12699
rect 17276 12668 17325 12696
rect 17276 12656 17282 12668
rect 17313 12665 17325 12668
rect 17359 12665 17371 12699
rect 21192 12696 21220 12724
rect 21358 12696 21364 12708
rect 21192 12668 21364 12696
rect 17313 12659 17371 12665
rect 21358 12656 21364 12668
rect 21416 12656 21422 12708
rect 20714 12628 20720 12640
rect 14476 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 21082 12588 21088 12640
rect 21140 12588 21146 12640
rect 22186 12588 22192 12640
rect 22244 12628 22250 12640
rect 22373 12631 22431 12637
rect 22373 12628 22385 12631
rect 22244 12600 22385 12628
rect 22244 12588 22250 12600
rect 22373 12597 22385 12600
rect 22419 12597 22431 12631
rect 22373 12591 22431 12597
rect 552 12538 23368 12560
rect 552 12486 19022 12538
rect 19074 12486 19086 12538
rect 19138 12486 19150 12538
rect 19202 12486 19214 12538
rect 19266 12486 19278 12538
rect 19330 12486 23368 12538
rect 552 12464 23368 12486
rect 4246 12384 4252 12436
rect 4304 12424 4310 12436
rect 4801 12427 4859 12433
rect 4801 12424 4813 12427
rect 4304 12396 4813 12424
rect 4304 12384 4310 12396
rect 4801 12393 4813 12396
rect 4847 12393 4859 12427
rect 4801 12387 4859 12393
rect 5258 12384 5264 12436
rect 5316 12384 5322 12436
rect 5902 12384 5908 12436
rect 5960 12384 5966 12436
rect 7466 12384 7472 12436
rect 7524 12384 7530 12436
rect 7834 12384 7840 12436
rect 7892 12384 7898 12436
rect 8386 12384 8392 12436
rect 8444 12424 8450 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8444 12396 8585 12424
rect 8444 12384 8450 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 8573 12387 8631 12393
rect 10778 12384 10784 12436
rect 10836 12384 10842 12436
rect 12894 12384 12900 12436
rect 12952 12384 12958 12436
rect 13633 12427 13691 12433
rect 13633 12393 13645 12427
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 5169 12359 5227 12365
rect 5169 12325 5181 12359
rect 5215 12356 5227 12359
rect 5534 12356 5540 12368
rect 5215 12328 5540 12356
rect 5215 12325 5227 12328
rect 5169 12319 5227 12325
rect 5534 12316 5540 12328
rect 5592 12356 5598 12368
rect 5920 12356 5948 12384
rect 7852 12356 7880 12384
rect 5592 12328 5948 12356
rect 7668 12328 7880 12356
rect 5592 12316 5598 12328
rect 7668 12297 7696 12328
rect 8478 12316 8484 12368
rect 8536 12316 8542 12368
rect 9668 12359 9726 12365
rect 9668 12325 9680 12359
rect 9714 12356 9726 12359
rect 9858 12356 9864 12368
rect 9714 12328 9864 12356
rect 9714 12325 9726 12328
rect 9668 12319 9726 12325
rect 9858 12316 9864 12328
rect 9916 12316 9922 12368
rect 9950 12316 9956 12368
rect 10008 12316 10014 12368
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 12078 12359 12136 12365
rect 12078 12356 12090 12359
rect 11572 12328 12090 12356
rect 11572 12316 11578 12328
rect 12078 12325 12090 12328
rect 12124 12325 12136 12359
rect 12078 12319 12136 12325
rect 12342 12316 12348 12368
rect 12400 12356 12406 12368
rect 12805 12359 12863 12365
rect 12805 12356 12817 12359
rect 12400 12328 12817 12356
rect 12400 12316 12406 12328
rect 12805 12325 12817 12328
rect 12851 12325 12863 12359
rect 13648 12356 13676 12387
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 14366 12424 14372 12436
rect 13780 12396 14372 12424
rect 13780 12384 13786 12396
rect 14366 12384 14372 12396
rect 14424 12384 14430 12436
rect 20346 12384 20352 12436
rect 20404 12424 20410 12436
rect 20993 12427 21051 12433
rect 20993 12424 21005 12427
rect 20404 12396 21005 12424
rect 20404 12384 20410 12396
rect 20993 12393 21005 12396
rect 21039 12424 21051 12427
rect 21821 12427 21879 12433
rect 21039 12396 21772 12424
rect 21039 12393 21051 12396
rect 20993 12387 21051 12393
rect 13970 12359 14028 12365
rect 13970 12356 13982 12359
rect 13648 12328 13982 12356
rect 12805 12319 12863 12325
rect 13970 12325 13982 12328
rect 14016 12325 14028 12359
rect 13970 12319 14028 12325
rect 16298 12316 16304 12368
rect 16356 12356 16362 12368
rect 17313 12359 17371 12365
rect 16356 12328 17264 12356
rect 16356 12316 16362 12328
rect 7653 12291 7711 12297
rect 7653 12257 7665 12291
rect 7699 12257 7711 12291
rect 7653 12251 7711 12257
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12257 7895 12291
rect 7837 12251 7895 12257
rect 5442 12180 5448 12232
rect 5500 12180 5506 12232
rect 7852 12152 7880 12251
rect 7926 12248 7932 12300
rect 7984 12248 7990 12300
rect 8496 12288 8524 12316
rect 8573 12291 8631 12297
rect 8573 12288 8585 12291
rect 8496 12260 8585 12288
rect 8573 12257 8585 12260
rect 8619 12257 8631 12291
rect 8573 12251 8631 12257
rect 8757 12291 8815 12297
rect 8757 12257 8769 12291
rect 8803 12288 8815 12291
rect 9968 12288 9996 12316
rect 17236 12300 17264 12328
rect 17313 12325 17325 12359
rect 17359 12356 17371 12359
rect 17359 12328 18184 12356
rect 17359 12325 17371 12328
rect 17313 12319 17371 12325
rect 8803 12260 9996 12288
rect 8803 12257 8815 12260
rect 8757 12251 8815 12257
rect 7944 12220 7972 12248
rect 8772 12220 8800 12251
rect 13446 12248 13452 12300
rect 13504 12248 13510 12300
rect 13814 12288 13820 12300
rect 13556 12260 13820 12288
rect 7944 12192 8800 12220
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12189 12403 12223
rect 12345 12183 12403 12189
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 13556 12220 13584 12260
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 15378 12248 15384 12300
rect 15436 12248 15442 12300
rect 16942 12248 16948 12300
rect 17000 12248 17006 12300
rect 17218 12248 17224 12300
rect 17276 12248 17282 12300
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12288 17463 12291
rect 17770 12288 17776 12300
rect 17451 12260 17776 12288
rect 17451 12257 17463 12260
rect 17405 12251 17463 12257
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 18156 12297 18184 12328
rect 21082 12316 21088 12368
rect 21140 12356 21146 12368
rect 21269 12359 21327 12365
rect 21269 12356 21281 12359
rect 21140 12328 21281 12356
rect 21140 12316 21146 12328
rect 21269 12325 21281 12328
rect 21315 12325 21327 12359
rect 21744 12356 21772 12396
rect 21821 12393 21833 12427
rect 21867 12424 21879 12427
rect 21910 12424 21916 12436
rect 21867 12396 21916 12424
rect 21867 12393 21879 12396
rect 21821 12387 21879 12393
rect 21910 12384 21916 12396
rect 21968 12424 21974 12436
rect 21968 12396 22600 12424
rect 21968 12384 21974 12396
rect 21744 12328 22416 12356
rect 21269 12319 21327 12325
rect 18141 12291 18199 12297
rect 18141 12257 18153 12291
rect 18187 12257 18199 12291
rect 18141 12251 18199 12257
rect 18325 12291 18383 12297
rect 18325 12257 18337 12291
rect 18371 12288 18383 12291
rect 18782 12288 18788 12300
rect 18371 12260 18788 12288
rect 18371 12257 18383 12260
rect 18325 12251 18383 12257
rect 18782 12248 18788 12260
rect 18840 12248 18846 12300
rect 20806 12248 20812 12300
rect 20864 12248 20870 12300
rect 20898 12248 20904 12300
rect 20956 12288 20962 12300
rect 21545 12291 21603 12297
rect 21545 12288 21557 12291
rect 20956 12260 21557 12288
rect 20956 12248 20962 12260
rect 21545 12257 21557 12260
rect 21591 12257 21603 12291
rect 21545 12251 21603 12257
rect 22005 12291 22063 12297
rect 22005 12257 22017 12291
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 22097 12291 22155 12297
rect 22097 12257 22109 12291
rect 22143 12288 22155 12291
rect 22186 12288 22192 12300
rect 22143 12260 22192 12288
rect 22143 12257 22155 12260
rect 22097 12251 22155 12257
rect 13127 12192 13584 12220
rect 13725 12223 13783 12229
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13725 12189 13737 12223
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 8202 12152 8208 12164
rect 7852 12124 8208 12152
rect 8202 12112 8208 12124
rect 8260 12112 8266 12164
rect 9416 12084 9444 12183
rect 12360 12152 12388 12183
rect 12360 12124 13676 12152
rect 13648 12096 13676 12124
rect 9582 12084 9588 12096
rect 9416 12056 9588 12084
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 10962 12044 10968 12096
rect 11020 12044 11026 12096
rect 12434 12044 12440 12096
rect 12492 12044 12498 12096
rect 13630 12044 13636 12096
rect 13688 12044 13694 12096
rect 13740 12084 13768 12183
rect 16850 12180 16856 12232
rect 16908 12220 16914 12232
rect 17083 12223 17141 12229
rect 17083 12220 17095 12223
rect 16908 12192 17095 12220
rect 16908 12180 16914 12192
rect 17083 12189 17095 12192
rect 17129 12220 17141 12223
rect 17678 12220 17684 12232
rect 17129 12192 17684 12220
rect 17129 12189 17141 12192
rect 17083 12183 17141 12189
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 20824 12152 20852 12248
rect 20990 12180 20996 12232
rect 21048 12220 21054 12232
rect 21361 12223 21419 12229
rect 21361 12220 21373 12223
rect 21048 12192 21373 12220
rect 21048 12180 21054 12192
rect 21361 12189 21373 12192
rect 21407 12189 21419 12223
rect 22020 12220 22048 12251
rect 22186 12248 22192 12260
rect 22244 12248 22250 12300
rect 22278 12248 22284 12300
rect 22336 12248 22342 12300
rect 21361 12183 21419 12189
rect 21744 12192 22048 12220
rect 22388 12220 22416 12328
rect 22572 12297 22600 12396
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12257 22615 12291
rect 22557 12251 22615 12257
rect 23017 12291 23075 12297
rect 23017 12257 23029 12291
rect 23063 12288 23075 12291
rect 23290 12288 23296 12300
rect 23063 12260 23296 12288
rect 23063 12257 23075 12260
rect 23017 12251 23075 12257
rect 23290 12248 23296 12260
rect 23348 12248 23354 12300
rect 22741 12223 22799 12229
rect 22741 12220 22753 12223
rect 22388 12192 22753 12220
rect 21744 12161 21772 12192
rect 22741 12189 22753 12192
rect 22787 12189 22799 12223
rect 22741 12183 22799 12189
rect 21729 12155 21787 12161
rect 20824 12124 21404 12152
rect 14366 12084 14372 12096
rect 13740 12056 14372 12084
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 15102 12044 15108 12096
rect 15160 12044 15166 12096
rect 15194 12044 15200 12096
rect 15252 12044 15258 12096
rect 18230 12044 18236 12096
rect 18288 12044 18294 12096
rect 21266 12044 21272 12096
rect 21324 12044 21330 12096
rect 21376 12084 21404 12124
rect 21729 12121 21741 12155
rect 21775 12121 21787 12155
rect 22833 12155 22891 12161
rect 22833 12152 22845 12155
rect 21729 12115 21787 12121
rect 21836 12124 22845 12152
rect 21836 12084 21864 12124
rect 22833 12121 22845 12124
rect 22879 12121 22891 12155
rect 22833 12115 22891 12121
rect 21376 12056 21864 12084
rect 22094 12044 22100 12096
rect 22152 12044 22158 12096
rect 22370 12044 22376 12096
rect 22428 12044 22434 12096
rect 552 11994 23368 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 23368 11994
rect 552 11920 23368 11942
rect 5353 11883 5411 11889
rect 5353 11849 5365 11883
rect 5399 11880 5411 11883
rect 5718 11880 5724 11892
rect 5399 11852 5724 11880
rect 5399 11849 5411 11852
rect 5353 11843 5411 11849
rect 5718 11840 5724 11852
rect 5776 11880 5782 11892
rect 5997 11883 6055 11889
rect 5997 11880 6009 11883
rect 5776 11852 6009 11880
rect 5776 11840 5782 11852
rect 5997 11849 6009 11852
rect 6043 11849 6055 11883
rect 5997 11843 6055 11849
rect 11054 11840 11060 11892
rect 11112 11880 11118 11892
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 11112 11852 11529 11880
rect 11112 11840 11118 11852
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 12434 11880 12440 11892
rect 11517 11843 11575 11849
rect 12406 11840 12440 11880
rect 12492 11840 12498 11892
rect 13541 11883 13599 11889
rect 13541 11849 13553 11883
rect 13587 11880 13599 11883
rect 13906 11880 13912 11892
rect 13587 11852 13912 11880
rect 13587 11849 13599 11852
rect 13541 11843 13599 11849
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 15102 11840 15108 11892
rect 15160 11840 15166 11892
rect 15194 11840 15200 11892
rect 15252 11840 15258 11892
rect 18230 11840 18236 11892
rect 18288 11840 18294 11892
rect 19245 11883 19303 11889
rect 19245 11849 19257 11883
rect 19291 11880 19303 11883
rect 19981 11883 20039 11889
rect 19981 11880 19993 11883
rect 19291 11852 19993 11880
rect 19291 11849 19303 11852
rect 19245 11843 19303 11849
rect 19981 11849 19993 11852
rect 20027 11849 20039 11883
rect 19981 11843 20039 11849
rect 20441 11883 20499 11889
rect 20441 11849 20453 11883
rect 20487 11880 20499 11883
rect 20898 11880 20904 11892
rect 20487 11852 20904 11880
rect 20487 11849 20499 11852
rect 20441 11843 20499 11849
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 20993 11883 21051 11889
rect 20993 11849 21005 11883
rect 21039 11880 21051 11883
rect 21450 11880 21456 11892
rect 21039 11852 21456 11880
rect 21039 11849 21051 11852
rect 20993 11843 21051 11849
rect 21450 11840 21456 11852
rect 21508 11840 21514 11892
rect 5534 11812 5540 11824
rect 5184 11784 5540 11812
rect 5184 11753 5212 11784
rect 5534 11772 5540 11784
rect 5592 11772 5598 11824
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5552 11744 5580 11772
rect 6089 11747 6147 11753
rect 6089 11744 6101 11747
rect 5552 11716 6101 11744
rect 5552 11685 5580 11716
rect 6089 11713 6101 11716
rect 6135 11713 6147 11747
rect 6089 11707 6147 11713
rect 10962 11704 10968 11756
rect 11020 11744 11026 11756
rect 11149 11747 11207 11753
rect 11149 11744 11161 11747
rect 11020 11716 11161 11744
rect 11020 11704 11026 11716
rect 11149 11713 11161 11716
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 5445 11679 5503 11685
rect 5445 11645 5457 11679
rect 5491 11645 5503 11679
rect 5445 11639 5503 11645
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11645 5595 11679
rect 5537 11639 5595 11645
rect 5460 11608 5488 11639
rect 5626 11636 5632 11688
rect 5684 11636 5690 11688
rect 5994 11636 6000 11688
rect 6052 11636 6058 11688
rect 6273 11679 6331 11685
rect 6273 11645 6285 11679
rect 6319 11645 6331 11679
rect 6273 11639 6331 11645
rect 5644 11608 5672 11636
rect 6288 11608 6316 11639
rect 6454 11636 6460 11688
rect 6512 11676 6518 11688
rect 7650 11676 7656 11688
rect 6512 11648 7656 11676
rect 6512 11636 6518 11648
rect 7650 11636 7656 11648
rect 7708 11676 7714 11688
rect 7929 11679 7987 11685
rect 7929 11676 7941 11679
rect 7708 11648 7941 11676
rect 7708 11636 7714 11648
rect 7929 11645 7941 11648
rect 7975 11645 7987 11679
rect 7929 11639 7987 11645
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11645 8171 11679
rect 8113 11639 8171 11645
rect 8128 11608 8156 11639
rect 11330 11636 11336 11688
rect 11388 11636 11394 11688
rect 12161 11679 12219 11685
rect 12161 11645 12173 11679
rect 12207 11676 12219 11679
rect 12406 11676 12434 11840
rect 15212 11812 15240 11840
rect 14936 11784 15240 11812
rect 15565 11815 15623 11821
rect 14936 11744 14964 11784
rect 15565 11781 15577 11815
rect 15611 11812 15623 11815
rect 16209 11815 16267 11821
rect 15611 11784 16068 11812
rect 15611 11781 15623 11784
rect 15565 11775 15623 11781
rect 14844 11716 14964 11744
rect 12207 11648 12434 11676
rect 14665 11679 14723 11685
rect 12207 11645 12219 11648
rect 12161 11639 12219 11645
rect 14665 11645 14677 11679
rect 14711 11676 14723 11679
rect 14844 11676 14872 11716
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15930 11744 15936 11756
rect 15344 11716 15936 11744
rect 15344 11704 15350 11716
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 16040 11744 16068 11784
rect 16209 11781 16221 11815
rect 16255 11812 16267 11815
rect 16255 11784 16436 11812
rect 16255 11781 16267 11784
rect 16209 11775 16267 11781
rect 16408 11756 16436 11784
rect 17218 11772 17224 11824
rect 17276 11772 17282 11824
rect 16298 11744 16304 11756
rect 16040 11716 16304 11744
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 16390 11704 16396 11756
rect 16448 11704 16454 11756
rect 17236 11744 17264 11772
rect 17144 11716 17264 11744
rect 18248 11744 18276 11840
rect 19889 11815 19947 11821
rect 19889 11781 19901 11815
rect 19935 11812 19947 11815
rect 19935 11784 20116 11812
rect 19935 11781 19947 11784
rect 19889 11775 19947 11781
rect 18785 11747 18843 11753
rect 18785 11744 18797 11747
rect 18248 11716 18797 11744
rect 14711 11648 14872 11676
rect 14921 11679 14979 11685
rect 14711 11645 14723 11648
rect 14665 11639 14723 11645
rect 14921 11645 14933 11679
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 15381 11679 15439 11685
rect 15381 11645 15393 11679
rect 15427 11645 15439 11679
rect 15381 11639 15439 11645
rect 16025 11679 16083 11685
rect 16025 11645 16037 11679
rect 16071 11645 16083 11679
rect 16025 11639 16083 11645
rect 16209 11679 16267 11685
rect 16209 11645 16221 11679
rect 16255 11676 16267 11679
rect 16316 11676 16344 11704
rect 16255 11648 16344 11676
rect 16563 11679 16621 11685
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 16563 11645 16575 11679
rect 16609 11676 16621 11679
rect 16850 11676 16856 11688
rect 16609 11648 16856 11676
rect 16609 11645 16621 11648
rect 16563 11639 16621 11645
rect 8570 11608 8576 11620
rect 5460 11580 6316 11608
rect 7208 11580 8576 11608
rect 7208 11552 7236 11580
rect 8570 11568 8576 11580
rect 8628 11568 8634 11620
rect 13814 11568 13820 11620
rect 13872 11608 13878 11620
rect 14936 11608 14964 11639
rect 13872 11580 14964 11608
rect 13872 11568 13878 11580
rect 14568 11552 14596 11580
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 15105 11611 15163 11617
rect 15105 11608 15117 11611
rect 15068 11580 15117 11608
rect 15068 11568 15074 11580
rect 15105 11577 15117 11580
rect 15151 11577 15163 11611
rect 15105 11571 15163 11577
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11540 5227 11543
rect 5810 11540 5816 11552
rect 5215 11512 5816 11540
rect 5215 11509 5227 11512
rect 5169 11503 5227 11509
rect 5810 11500 5816 11512
rect 5868 11500 5874 11552
rect 5902 11500 5908 11552
rect 5960 11500 5966 11552
rect 6457 11543 6515 11549
rect 6457 11509 6469 11543
rect 6503 11540 6515 11543
rect 7190 11540 7196 11552
rect 6503 11512 7196 11540
rect 6503 11509 6515 11512
rect 6457 11503 6515 11509
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 8021 11543 8079 11549
rect 8021 11509 8033 11543
rect 8067 11540 8079 11543
rect 8662 11540 8668 11552
rect 8067 11512 8668 11540
rect 8067 11509 8079 11512
rect 8021 11503 8079 11509
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 11974 11500 11980 11552
rect 12032 11500 12038 11552
rect 14550 11500 14556 11552
rect 14608 11500 14614 11552
rect 14734 11500 14740 11552
rect 14792 11540 14798 11552
rect 15396 11540 15424 11639
rect 16040 11608 16068 11639
rect 16850 11636 16856 11648
rect 16908 11636 16914 11688
rect 16942 11636 16948 11688
rect 17000 11636 17006 11688
rect 17144 11687 17172 11716
rect 18785 11713 18797 11716
rect 18831 11713 18843 11747
rect 18785 11707 18843 11713
rect 19426 11704 19432 11756
rect 19484 11704 19490 11756
rect 20088 11753 20116 11784
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11713 20131 11747
rect 20073 11707 20131 11713
rect 17129 11681 17187 11687
rect 17129 11647 17141 11681
rect 17175 11647 17187 11681
rect 17129 11641 17187 11647
rect 17221 11679 17279 11685
rect 17221 11645 17233 11679
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11645 18935 11679
rect 18877 11639 18935 11645
rect 16960 11608 16988 11636
rect 17236 11608 17264 11639
rect 16040 11580 17264 11608
rect 18782 11568 18788 11620
rect 18840 11608 18846 11620
rect 18892 11608 18920 11639
rect 19518 11636 19524 11688
rect 19576 11636 19582 11688
rect 20254 11636 20260 11688
rect 20312 11636 20318 11688
rect 22373 11679 22431 11685
rect 22373 11645 22385 11679
rect 22419 11676 22431 11679
rect 22554 11676 22560 11688
rect 22419 11648 22560 11676
rect 22419 11645 22431 11648
rect 22373 11639 22431 11645
rect 22554 11636 22560 11648
rect 22612 11636 22618 11688
rect 18840 11580 18920 11608
rect 18840 11568 18846 11580
rect 19978 11568 19984 11620
rect 20036 11568 20042 11620
rect 22128 11611 22186 11617
rect 22128 11577 22140 11611
rect 22174 11608 22186 11611
rect 22278 11608 22284 11620
rect 22174 11580 22284 11608
rect 22174 11577 22186 11580
rect 22128 11571 22186 11577
rect 22278 11568 22284 11580
rect 22336 11568 22342 11620
rect 14792 11512 15424 11540
rect 14792 11500 14798 11512
rect 16850 11500 16856 11552
rect 16908 11500 16914 11552
rect 16942 11500 16948 11552
rect 17000 11500 17006 11552
rect 20990 11500 20996 11552
rect 21048 11540 21054 11552
rect 22370 11540 22376 11552
rect 21048 11512 22376 11540
rect 21048 11500 21054 11512
rect 22370 11500 22376 11512
rect 22428 11500 22434 11552
rect 552 11450 23368 11472
rect 552 11398 19022 11450
rect 19074 11398 19086 11450
rect 19138 11398 19150 11450
rect 19202 11398 19214 11450
rect 19266 11398 19278 11450
rect 19330 11398 23368 11450
rect 552 11376 23368 11398
rect 6178 11296 6184 11348
rect 6236 11336 6242 11348
rect 6825 11339 6883 11345
rect 6236 11308 6592 11336
rect 6236 11296 6242 11308
rect 5442 11228 5448 11280
rect 5500 11268 5506 11280
rect 6564 11277 6592 11308
rect 6825 11305 6837 11339
rect 6871 11336 6883 11339
rect 7282 11336 7288 11348
rect 7340 11345 7346 11348
rect 7340 11339 7359 11345
rect 6871 11308 7288 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 7282 11296 7288 11308
rect 7347 11305 7359 11339
rect 7340 11299 7359 11305
rect 9033 11339 9091 11345
rect 9033 11305 9045 11339
rect 9079 11336 9091 11339
rect 9674 11336 9680 11348
rect 9079 11308 9680 11336
rect 9079 11305 9091 11308
rect 9033 11299 9091 11305
rect 7340 11296 7346 11299
rect 9674 11296 9680 11308
rect 9732 11336 9738 11348
rect 9732 11308 11284 11336
rect 9732 11296 9738 11308
rect 5813 11271 5871 11277
rect 5813 11268 5825 11271
rect 5500 11240 5825 11268
rect 5500 11228 5506 11240
rect 5813 11237 5825 11240
rect 5859 11237 5871 11271
rect 5813 11231 5871 11237
rect 6029 11271 6087 11277
rect 6029 11237 6041 11271
rect 6075 11268 6087 11271
rect 6549 11271 6607 11277
rect 6075 11240 6224 11268
rect 6075 11237 6087 11240
rect 6029 11231 6087 11237
rect 5261 11203 5319 11209
rect 5261 11169 5273 11203
rect 5307 11200 5319 11203
rect 5718 11200 5724 11212
rect 5307 11172 5724 11200
rect 5307 11169 5319 11172
rect 5261 11163 5319 11169
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 6196 11200 6224 11240
rect 6549 11237 6561 11271
rect 6595 11237 6607 11271
rect 6549 11231 6607 11237
rect 7101 11271 7159 11277
rect 7101 11237 7113 11271
rect 7147 11268 7159 11271
rect 7558 11268 7564 11280
rect 7147 11240 7564 11268
rect 7147 11237 7159 11240
rect 7101 11231 7159 11237
rect 7558 11228 7564 11240
rect 7616 11228 7622 11280
rect 7668 11240 8432 11268
rect 7668 11212 7696 11240
rect 6273 11203 6331 11209
rect 6273 11200 6285 11203
rect 5828 11172 6285 11200
rect 5828 11144 5856 11172
rect 6273 11169 6285 11172
rect 6319 11169 6331 11203
rect 6273 11163 6331 11169
rect 6365 11203 6423 11209
rect 6365 11169 6377 11203
rect 6411 11169 6423 11203
rect 6365 11163 6423 11169
rect 6641 11203 6699 11209
rect 6641 11169 6653 11203
rect 6687 11169 6699 11203
rect 6641 11163 6699 11169
rect 6825 11203 6883 11209
rect 6825 11169 6837 11203
rect 6871 11169 6883 11203
rect 6825 11163 6883 11169
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 5368 11064 5396 11095
rect 5810 11092 5816 11144
rect 5868 11092 5874 11144
rect 6380 11132 6408 11163
rect 6656 11132 6684 11163
rect 6012 11104 6684 11132
rect 5718 11064 5724 11076
rect 5368 11036 5724 11064
rect 5718 11024 5724 11036
rect 5776 11024 5782 11076
rect 5534 10956 5540 11008
rect 5592 10956 5598 11008
rect 5902 10956 5908 11008
rect 5960 10996 5966 11008
rect 6012 11005 6040 11104
rect 6086 11024 6092 11076
rect 6144 11064 6150 11076
rect 6840 11064 6868 11163
rect 7650 11160 7656 11212
rect 7708 11160 7714 11212
rect 8036 11209 8064 11240
rect 8202 11209 8208 11212
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 8159 11203 8208 11209
rect 8159 11169 8171 11203
rect 8205 11169 8208 11203
rect 8159 11163 8208 11169
rect 7760 11132 7788 11163
rect 8202 11160 8208 11163
rect 8260 11160 8266 11212
rect 8297 11135 8355 11141
rect 8297 11132 8309 11135
rect 6144 11036 6868 11064
rect 7300 11104 8309 11132
rect 6144 11024 6150 11036
rect 5997 10999 6055 11005
rect 5997 10996 6009 10999
rect 5960 10968 6009 10996
rect 5960 10956 5966 10968
rect 5997 10965 6009 10968
rect 6043 10965 6055 10999
rect 5997 10959 6055 10965
rect 6181 10999 6239 11005
rect 6181 10965 6193 10999
rect 6227 10996 6239 10999
rect 6270 10996 6276 11008
rect 6227 10968 6276 10996
rect 6227 10965 6239 10968
rect 6181 10959 6239 10965
rect 6270 10956 6276 10968
rect 6328 10956 6334 11008
rect 6546 10956 6552 11008
rect 6604 10956 6610 11008
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 7300 11005 7328 11104
rect 8297 11101 8309 11104
rect 8343 11101 8355 11135
rect 8404 11132 8432 11240
rect 8570 11228 8576 11280
rect 8628 11228 8634 11280
rect 8478 11160 8484 11212
rect 8536 11200 8542 11212
rect 8757 11203 8815 11209
rect 8757 11200 8769 11203
rect 8536 11172 8769 11200
rect 8536 11160 8542 11172
rect 8757 11169 8769 11172
rect 8803 11169 8815 11203
rect 8757 11163 8815 11169
rect 8849 11203 8907 11209
rect 8849 11169 8861 11203
rect 8895 11169 8907 11203
rect 8849 11163 8907 11169
rect 8864 11132 8892 11163
rect 10778 11160 10784 11212
rect 10836 11200 10842 11212
rect 11256 11209 11284 11308
rect 11974 11296 11980 11348
rect 12032 11296 12038 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 12897 11339 12955 11345
rect 12897 11336 12909 11339
rect 12400 11308 12909 11336
rect 12400 11296 12406 11308
rect 12897 11305 12909 11308
rect 12943 11305 12955 11339
rect 12897 11299 12955 11305
rect 16298 11296 16304 11348
rect 16356 11296 16362 11348
rect 16942 11296 16948 11348
rect 17000 11296 17006 11348
rect 19978 11296 19984 11348
rect 20036 11296 20042 11348
rect 20901 11339 20959 11345
rect 20901 11305 20913 11339
rect 20947 11336 20959 11339
rect 20990 11336 20996 11348
rect 20947 11308 20996 11336
rect 20947 11305 20959 11308
rect 20901 11299 20959 11305
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 21085 11339 21143 11345
rect 21085 11305 21097 11339
rect 21131 11336 21143 11339
rect 22094 11336 22100 11348
rect 21131 11308 22100 11336
rect 21131 11305 21143 11308
rect 21085 11299 21143 11305
rect 22094 11296 22100 11308
rect 22152 11296 22158 11348
rect 22649 11339 22707 11345
rect 22649 11305 22661 11339
rect 22695 11305 22707 11339
rect 22649 11299 22707 11305
rect 11784 11271 11842 11277
rect 11348 11240 11744 11268
rect 11348 11209 11376 11240
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 10836 11172 10977 11200
rect 10836 11160 10842 11172
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11241 11203 11299 11209
rect 11241 11169 11253 11203
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11169 11483 11203
rect 11716 11200 11744 11240
rect 11784 11237 11796 11271
rect 11830 11268 11842 11271
rect 11992 11268 12020 11296
rect 15105 11271 15163 11277
rect 11830 11240 12020 11268
rect 14016 11240 14320 11268
rect 11830 11237 11842 11240
rect 11784 11231 11842 11237
rect 12618 11200 12624 11212
rect 11716 11172 12624 11200
rect 11425 11163 11483 11169
rect 8404 11104 8892 11132
rect 8297 11095 8355 11101
rect 7929 11067 7987 11073
rect 7929 11033 7941 11067
rect 7975 11064 7987 11067
rect 9858 11064 9864 11076
rect 7975 11036 9864 11064
rect 7975 11033 7987 11036
rect 7929 11027 7987 11033
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 10962 11024 10968 11076
rect 11020 11064 11026 11076
rect 11103 11067 11161 11073
rect 11103 11064 11115 11067
rect 11020 11036 11115 11064
rect 11020 11024 11026 11036
rect 11103 11033 11115 11036
rect 11149 11033 11161 11067
rect 11103 11027 11161 11033
rect 7285 10999 7343 11005
rect 7285 10996 7297 10999
rect 7248 10968 7297 10996
rect 7248 10956 7254 10968
rect 7285 10965 7297 10968
rect 7331 10965 7343 10999
rect 7285 10959 7343 10965
rect 7469 10999 7527 11005
rect 7469 10965 7481 10999
rect 7515 10996 7527 10999
rect 7834 10996 7840 11008
rect 7515 10968 7840 10996
rect 7515 10965 7527 10968
rect 7469 10959 7527 10965
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 8386 10956 8392 11008
rect 8444 10956 8450 11008
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 8573 10999 8631 11005
rect 8573 10996 8585 10999
rect 8536 10968 8585 10996
rect 8536 10956 8542 10968
rect 8573 10965 8585 10968
rect 8619 10965 8631 10999
rect 8573 10959 8631 10965
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 10042 10996 10048 11008
rect 8720 10968 10048 10996
rect 8720 10956 8726 10968
rect 10042 10956 10048 10968
rect 10100 10956 10106 11008
rect 11440 10996 11468 11163
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 13906 11160 13912 11212
rect 13964 11200 13970 11212
rect 14016 11209 14044 11240
rect 14292 11212 14320 11240
rect 15105 11237 15117 11271
rect 15151 11268 15163 11271
rect 15151 11240 16160 11268
rect 15151 11237 15163 11240
rect 15105 11231 15163 11237
rect 14001 11203 14059 11209
rect 14001 11200 14013 11203
rect 13964 11172 14013 11200
rect 13964 11160 13970 11172
rect 14001 11169 14013 11172
rect 14047 11169 14059 11203
rect 14001 11163 14059 11169
rect 14090 11160 14096 11212
rect 14148 11200 14154 11212
rect 14185 11203 14243 11209
rect 14185 11200 14197 11203
rect 14148 11172 14197 11200
rect 14148 11160 14154 11172
rect 14185 11169 14197 11172
rect 14231 11169 14243 11203
rect 14185 11163 14243 11169
rect 11514 11092 11520 11144
rect 11572 11092 11578 11144
rect 14200 11132 14228 11163
rect 14274 11160 14280 11212
rect 14332 11200 14338 11212
rect 14734 11200 14740 11212
rect 14332 11172 14740 11200
rect 14332 11160 14338 11172
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 15197 11203 15255 11209
rect 15197 11169 15209 11203
rect 15243 11200 15255 11203
rect 15286 11200 15292 11212
rect 15243 11172 15292 11200
rect 15243 11169 15255 11172
rect 15197 11163 15255 11169
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 16132 11209 16160 11240
rect 16316 11209 16344 11296
rect 16117 11203 16175 11209
rect 16117 11169 16129 11203
rect 16163 11169 16175 11203
rect 16117 11163 16175 11169
rect 16301 11203 16359 11209
rect 16301 11169 16313 11203
rect 16347 11169 16359 11203
rect 16301 11163 16359 11169
rect 16390 11160 16396 11212
rect 16448 11200 16454 11212
rect 16577 11203 16635 11209
rect 16577 11200 16589 11203
rect 16448 11172 16589 11200
rect 16448 11160 16454 11172
rect 16577 11169 16589 11172
rect 16623 11169 16635 11203
rect 16577 11163 16635 11169
rect 16761 11203 16819 11209
rect 16761 11169 16773 11203
rect 16807 11200 16819 11203
rect 16960 11200 16988 11296
rect 16807 11172 16988 11200
rect 16807 11169 16819 11172
rect 16761 11163 16819 11169
rect 18874 11160 18880 11212
rect 18932 11160 18938 11212
rect 19886 11200 19892 11212
rect 18984 11172 19892 11200
rect 15010 11132 15016 11144
rect 14200 11104 15016 11132
rect 15010 11092 15016 11104
rect 15068 11092 15074 11144
rect 18984 11141 19012 11172
rect 19886 11160 19892 11172
rect 19944 11160 19950 11212
rect 18969 11135 19027 11141
rect 18969 11101 18981 11135
rect 19015 11101 19027 11135
rect 18969 11095 19027 11101
rect 19245 11135 19303 11141
rect 19245 11101 19257 11135
rect 19291 11132 19303 11135
rect 19996 11132 20024 11296
rect 21358 11228 21364 11280
rect 21416 11268 21422 11280
rect 22002 11268 22008 11280
rect 21416 11240 22008 11268
rect 21416 11228 21422 11240
rect 22002 11228 22008 11240
rect 22060 11268 22066 11280
rect 22664 11268 22692 11299
rect 22060 11240 22692 11268
rect 22060 11228 22066 11240
rect 21525 11203 21583 11209
rect 21525 11200 21537 11203
rect 20916 11172 21537 11200
rect 20916 11144 20944 11172
rect 21525 11169 21537 11172
rect 21571 11169 21583 11203
rect 21525 11163 21583 11169
rect 19291 11104 20024 11132
rect 19291 11101 19303 11104
rect 19245 11095 19303 11101
rect 20898 11092 20904 11144
rect 20956 11092 20962 11144
rect 21269 11135 21327 11141
rect 21269 11101 21281 11135
rect 21315 11101 21327 11135
rect 21269 11095 21327 11101
rect 14875 11067 14933 11073
rect 14875 11064 14887 11067
rect 14016 11036 14887 11064
rect 14016 11008 14044 11036
rect 14875 11033 14887 11036
rect 14921 11064 14933 11067
rect 15102 11064 15108 11076
rect 14921 11036 15108 11064
rect 14921 11033 14933 11036
rect 14875 11027 14933 11033
rect 15102 11024 15108 11036
rect 15160 11024 15166 11076
rect 20530 11024 20536 11076
rect 20588 11024 20594 11076
rect 21284 11064 21312 11095
rect 20824 11036 21312 11064
rect 11882 10996 11888 11008
rect 11440 10968 11888 10996
rect 11882 10956 11888 10968
rect 11940 10996 11946 11008
rect 12250 10996 12256 11008
rect 11940 10968 12256 10996
rect 11940 10956 11946 10968
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 13998 10956 14004 11008
rect 14056 10956 14062 11008
rect 14182 10956 14188 11008
rect 14240 10956 14246 11008
rect 16206 10956 16212 11008
rect 16264 10956 16270 11008
rect 16758 10956 16764 11008
rect 16816 10956 16822 11008
rect 19610 10956 19616 11008
rect 19668 10996 19674 11008
rect 20824 10996 20852 11036
rect 19668 10968 20852 10996
rect 20901 10999 20959 11005
rect 19668 10956 19674 10968
rect 20901 10965 20913 10999
rect 20947 10996 20959 10999
rect 20990 10996 20996 11008
rect 20947 10968 20996 10996
rect 20947 10965 20959 10968
rect 20901 10959 20959 10965
rect 20990 10956 20996 10968
rect 21048 10956 21054 11008
rect 552 10906 23368 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 23368 10906
rect 552 10832 23368 10854
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 6178 10792 6184 10804
rect 5500 10764 6184 10792
rect 5500 10752 5506 10764
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 6270 10752 6276 10804
rect 6328 10752 6334 10804
rect 8205 10795 8263 10801
rect 8205 10761 8217 10795
rect 8251 10792 8263 10795
rect 9033 10795 9091 10801
rect 9033 10792 9045 10795
rect 8251 10764 9045 10792
rect 8251 10761 8263 10764
rect 8205 10755 8263 10761
rect 9033 10761 9045 10764
rect 9079 10761 9091 10795
rect 9033 10755 9091 10761
rect 9674 10752 9680 10804
rect 9732 10752 9738 10804
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11020 10764 11713 10792
rect 11020 10752 11026 10764
rect 11701 10761 11713 10764
rect 11747 10761 11759 10795
rect 11701 10755 11759 10761
rect 16393 10795 16451 10801
rect 16393 10761 16405 10795
rect 16439 10792 16451 10795
rect 17773 10795 17831 10801
rect 17773 10792 17785 10795
rect 16439 10764 17785 10792
rect 16439 10761 16451 10764
rect 16393 10755 16451 10761
rect 17773 10761 17785 10764
rect 17819 10761 17831 10795
rect 17773 10755 17831 10761
rect 18233 10795 18291 10801
rect 18233 10761 18245 10795
rect 18279 10792 18291 10795
rect 20254 10792 20260 10804
rect 18279 10764 20260 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 20254 10752 20260 10764
rect 20312 10752 20318 10804
rect 20530 10752 20536 10804
rect 20588 10752 20594 10804
rect 20898 10752 20904 10804
rect 20956 10752 20962 10804
rect 20990 10752 20996 10804
rect 21048 10792 21054 10804
rect 21085 10795 21143 10801
rect 21085 10792 21097 10795
rect 21048 10764 21097 10792
rect 21048 10752 21054 10764
rect 21085 10761 21097 10764
rect 21131 10761 21143 10795
rect 21085 10755 21143 10761
rect 21821 10795 21879 10801
rect 21821 10761 21833 10795
rect 21867 10761 21879 10795
rect 21821 10755 21879 10761
rect 7745 10727 7803 10733
rect 7745 10693 7757 10727
rect 7791 10693 7803 10727
rect 7745 10687 7803 10693
rect 5534 10616 5540 10668
rect 5592 10616 5598 10668
rect 6546 10616 6552 10668
rect 6604 10616 6610 10668
rect 6638 10548 6644 10600
rect 6696 10548 6702 10600
rect 7282 10548 7288 10600
rect 7340 10588 7346 10600
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 7340 10560 7481 10588
rect 7340 10548 7346 10560
rect 7469 10557 7481 10560
rect 7515 10557 7527 10591
rect 7760 10588 7788 10687
rect 7834 10684 7840 10736
rect 7892 10684 7898 10736
rect 8386 10684 8392 10736
rect 8444 10724 8450 10736
rect 8444 10696 9628 10724
rect 8444 10684 8450 10696
rect 7852 10656 7880 10684
rect 7852 10628 8064 10656
rect 8036 10597 8064 10628
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 8260 10628 8616 10656
rect 8260 10616 8266 10628
rect 7837 10591 7895 10597
rect 7837 10588 7849 10591
rect 7760 10560 7849 10588
rect 7469 10551 7527 10557
rect 7837 10557 7849 10560
rect 7883 10557 7895 10591
rect 7837 10551 7895 10557
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10557 8079 10591
rect 8588 10588 8616 10628
rect 8662 10616 8668 10668
rect 8720 10616 8726 10668
rect 8864 10628 9352 10656
rect 8757 10591 8815 10597
rect 8757 10588 8769 10591
rect 8588 10560 8769 10588
rect 8021 10551 8079 10557
rect 8757 10557 8769 10560
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 5721 10523 5779 10529
rect 5721 10520 5733 10523
rect 5552 10492 5733 10520
rect 5552 10464 5580 10492
rect 5721 10489 5733 10492
rect 5767 10489 5779 10523
rect 6181 10523 6239 10529
rect 6181 10520 6193 10523
rect 5721 10483 5779 10489
rect 6104 10492 6193 10520
rect 5534 10412 5540 10464
rect 5592 10412 5598 10464
rect 5626 10412 5632 10464
rect 5684 10412 5690 10464
rect 6104 10461 6132 10492
rect 6181 10489 6193 10492
rect 6227 10489 6239 10523
rect 6181 10483 6239 10489
rect 6840 10492 7696 10520
rect 6840 10461 6868 10492
rect 6089 10455 6147 10461
rect 6089 10421 6101 10455
rect 6135 10421 6147 10455
rect 6089 10415 6147 10421
rect 6825 10455 6883 10461
rect 6825 10421 6837 10455
rect 6871 10421 6883 10455
rect 6825 10415 6883 10421
rect 7190 10412 7196 10464
rect 7248 10452 7254 10464
rect 7561 10455 7619 10461
rect 7561 10452 7573 10455
rect 7248 10424 7573 10452
rect 7248 10412 7254 10424
rect 7561 10421 7573 10424
rect 7607 10421 7619 10455
rect 7668 10452 7696 10492
rect 7742 10480 7748 10532
rect 7800 10480 7806 10532
rect 8864 10520 8892 10628
rect 9324 10597 9352 10628
rect 9600 10597 9628 10696
rect 9692 10656 9720 10752
rect 10594 10684 10600 10736
rect 10652 10724 10658 10736
rect 12161 10727 12219 10733
rect 10652 10696 11652 10724
rect 10652 10684 10658 10696
rect 10413 10659 10471 10665
rect 9692 10628 10364 10656
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10557 9275 10591
rect 9217 10551 9275 10557
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 9692 10588 9720 10628
rect 9769 10591 9827 10597
rect 9769 10588 9781 10591
rect 9692 10560 9781 10588
rect 9585 10551 9643 10557
rect 9769 10557 9781 10560
rect 9815 10557 9827 10591
rect 9769 10551 9827 10557
rect 8312 10492 8892 10520
rect 8312 10452 8340 10492
rect 9030 10480 9036 10532
rect 9088 10480 9094 10532
rect 9232 10520 9260 10551
rect 9858 10548 9864 10600
rect 9916 10548 9922 10600
rect 10042 10548 10048 10600
rect 10100 10548 10106 10600
rect 10336 10597 10364 10628
rect 10413 10625 10425 10659
rect 10459 10656 10471 10659
rect 10686 10656 10692 10668
rect 10459 10628 10692 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 10686 10616 10692 10628
rect 10744 10616 10750 10668
rect 11624 10665 11652 10696
rect 12161 10693 12173 10727
rect 12207 10724 12219 10727
rect 17037 10727 17095 10733
rect 12207 10696 12434 10724
rect 12207 10693 12219 10696
rect 12161 10687 12219 10693
rect 11609 10659 11667 10665
rect 11609 10625 11621 10659
rect 11655 10625 11667 10659
rect 11609 10619 11667 10625
rect 10321 10591 10379 10597
rect 10321 10557 10333 10591
rect 10367 10557 10379 10591
rect 10321 10551 10379 10557
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10588 10563 10591
rect 10594 10588 10600 10600
rect 10551 10560 10600 10588
rect 10551 10557 10563 10560
rect 10505 10551 10563 10557
rect 9232 10492 9444 10520
rect 9416 10464 9444 10492
rect 9674 10480 9680 10532
rect 9732 10520 9738 10532
rect 9953 10523 10011 10529
rect 9953 10520 9965 10523
rect 9732 10492 9965 10520
rect 9732 10480 9738 10492
rect 9953 10489 9965 10492
rect 9999 10489 10011 10523
rect 10336 10520 10364 10551
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10588 10839 10591
rect 10962 10588 10968 10600
rect 10827 10560 10968 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11425 10591 11483 10597
rect 11425 10557 11437 10591
rect 11471 10557 11483 10591
rect 11624 10588 11652 10619
rect 11882 10616 11888 10668
rect 11940 10616 11946 10668
rect 12406 10656 12434 10696
rect 17037 10693 17049 10727
rect 17083 10724 17095 10727
rect 20548 10724 20576 10752
rect 20714 10724 20720 10736
rect 17083 10696 17908 10724
rect 20548 10696 20720 10724
rect 17083 10693 17095 10696
rect 17037 10687 17095 10693
rect 14093 10659 14151 10665
rect 12406 10628 12848 10656
rect 11977 10591 12035 10597
rect 11977 10588 11989 10591
rect 11624 10560 11989 10588
rect 11425 10551 11483 10557
rect 11977 10557 11989 10560
rect 12023 10557 12035 10591
rect 11977 10551 12035 10557
rect 11440 10520 11468 10551
rect 12618 10548 12624 10600
rect 12676 10548 12682 10600
rect 12820 10597 12848 10628
rect 14093 10625 14105 10659
rect 14139 10656 14151 10659
rect 14182 10656 14188 10668
rect 14139 10628 14188 10656
rect 14139 10625 14151 10628
rect 14093 10619 14151 10625
rect 14182 10616 14188 10628
rect 14240 10656 14246 10668
rect 16117 10659 16175 10665
rect 14240 10628 14964 10656
rect 14240 10616 14246 10628
rect 12805 10591 12863 10597
rect 12805 10557 12817 10591
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 11701 10523 11759 10529
rect 11701 10520 11713 10523
rect 10336 10492 11713 10520
rect 9953 10483 10011 10489
rect 11701 10489 11713 10492
rect 11747 10489 11759 10523
rect 12820 10520 12848 10551
rect 13998 10548 14004 10600
rect 14056 10548 14062 10600
rect 14274 10548 14280 10600
rect 14332 10548 14338 10600
rect 14936 10597 14964 10628
rect 16117 10625 16129 10659
rect 16163 10656 16175 10659
rect 16206 10656 16212 10668
rect 16163 10628 16212 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 16758 10616 16764 10668
rect 16816 10616 16822 10668
rect 16850 10616 16856 10668
rect 16908 10656 16914 10668
rect 17880 10665 17908 10696
rect 20714 10684 20720 10696
rect 20772 10724 20778 10736
rect 21542 10724 21548 10736
rect 20772 10696 21548 10724
rect 20772 10684 20778 10696
rect 21542 10684 21548 10696
rect 21600 10724 21606 10736
rect 21637 10727 21695 10733
rect 21637 10724 21649 10727
rect 21600 10696 21649 10724
rect 21600 10684 21606 10696
rect 21637 10693 21649 10696
rect 21683 10693 21695 10727
rect 21637 10687 21695 10693
rect 17221 10659 17279 10665
rect 17221 10656 17233 10659
rect 16908 10628 17233 10656
rect 16908 10616 16914 10628
rect 17221 10625 17233 10628
rect 17267 10625 17279 10659
rect 17221 10619 17279 10625
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10625 17923 10659
rect 21836 10656 21864 10755
rect 22278 10752 22284 10804
rect 22336 10752 22342 10804
rect 17865 10619 17923 10625
rect 21468 10628 21864 10656
rect 21468 10600 21496 10628
rect 14461 10591 14519 10597
rect 14461 10557 14473 10591
rect 14507 10557 14519 10591
rect 14461 10551 14519 10557
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10588 14703 10591
rect 14737 10591 14795 10597
rect 14737 10588 14749 10591
rect 14691 10560 14749 10588
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 14737 10557 14749 10560
rect 14783 10557 14795 10591
rect 14737 10551 14795 10557
rect 14921 10591 14979 10597
rect 14921 10557 14933 10591
rect 14967 10557 14979 10591
rect 14921 10551 14979 10557
rect 14090 10520 14096 10532
rect 12820 10492 14096 10520
rect 11701 10483 11759 10489
rect 14090 10480 14096 10492
rect 14148 10520 14154 10532
rect 14476 10520 14504 10551
rect 16022 10548 16028 10600
rect 16080 10548 16086 10600
rect 16666 10548 16672 10600
rect 16724 10548 16730 10600
rect 17310 10548 17316 10600
rect 17368 10548 17374 10600
rect 18046 10548 18052 10600
rect 18104 10548 18110 10600
rect 20625 10591 20683 10597
rect 20625 10557 20637 10591
rect 20671 10588 20683 10591
rect 21269 10591 21327 10597
rect 20671 10560 21220 10588
rect 20671 10557 20683 10560
rect 20625 10551 20683 10557
rect 17773 10523 17831 10529
rect 17773 10520 17785 10523
rect 14148 10492 14504 10520
rect 17696 10492 17785 10520
rect 14148 10480 14154 10492
rect 7668 10424 8340 10452
rect 7561 10415 7619 10421
rect 8386 10412 8392 10464
rect 8444 10412 8450 10464
rect 9398 10412 9404 10464
rect 9456 10412 9462 10464
rect 9490 10412 9496 10464
rect 9548 10412 9554 10464
rect 9766 10412 9772 10464
rect 9824 10412 9830 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 11112 10424 11161 10452
rect 11112 10412 11118 10424
rect 11149 10421 11161 10424
rect 11195 10421 11207 10455
rect 11149 10415 11207 10421
rect 11238 10412 11244 10464
rect 11296 10412 11302 10464
rect 12802 10412 12808 10464
rect 12860 10412 12866 10464
rect 13633 10455 13691 10461
rect 13633 10421 13645 10455
rect 13679 10452 13691 10455
rect 13906 10452 13912 10464
rect 13679 10424 13912 10452
rect 13679 10421 13691 10424
rect 13633 10415 13691 10421
rect 13906 10412 13912 10424
rect 13964 10412 13970 10464
rect 14826 10412 14832 10464
rect 14884 10412 14890 10464
rect 17696 10461 17724 10492
rect 17773 10489 17785 10492
rect 17819 10489 17831 10523
rect 17773 10483 17831 10489
rect 20640 10464 20668 10551
rect 20898 10480 20904 10532
rect 20956 10480 20962 10532
rect 21192 10520 21220 10560
rect 21269 10557 21281 10591
rect 21315 10588 21327 10591
rect 21450 10588 21456 10600
rect 21315 10560 21456 10588
rect 21315 10557 21327 10560
rect 21269 10551 21327 10557
rect 21450 10548 21456 10560
rect 21508 10548 21514 10600
rect 21545 10591 21603 10597
rect 21545 10557 21557 10591
rect 21591 10557 21603 10591
rect 21545 10551 21603 10557
rect 21560 10520 21588 10551
rect 22094 10548 22100 10600
rect 22152 10548 22158 10600
rect 21789 10523 21847 10529
rect 21789 10520 21801 10523
rect 21192 10492 21801 10520
rect 21789 10489 21801 10492
rect 21835 10489 21847 10523
rect 21789 10483 21847 10489
rect 22002 10480 22008 10532
rect 22060 10480 22066 10532
rect 17681 10455 17739 10461
rect 17681 10421 17693 10455
rect 17727 10421 17739 10455
rect 17681 10415 17739 10421
rect 20622 10412 20628 10464
rect 20680 10412 20686 10464
rect 20717 10455 20775 10461
rect 20717 10421 20729 10455
rect 20763 10452 20775 10455
rect 21358 10452 21364 10464
rect 20763 10424 21364 10452
rect 20763 10421 20775 10424
rect 20717 10415 20775 10421
rect 21358 10412 21364 10424
rect 21416 10452 21422 10464
rect 21453 10455 21511 10461
rect 21453 10452 21465 10455
rect 21416 10424 21465 10452
rect 21416 10412 21422 10424
rect 21453 10421 21465 10424
rect 21499 10421 21511 10455
rect 21453 10415 21511 10421
rect 552 10362 23368 10384
rect 552 10310 19022 10362
rect 19074 10310 19086 10362
rect 19138 10310 19150 10362
rect 19202 10310 19214 10362
rect 19266 10310 19278 10362
rect 19330 10310 23368 10362
rect 552 10288 23368 10310
rect 6457 10251 6515 10257
rect 6457 10217 6469 10251
rect 6503 10248 6515 10251
rect 6638 10248 6644 10260
rect 6503 10220 6644 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 8386 10248 8392 10260
rect 8312 10220 8392 10248
rect 5258 10140 5264 10192
rect 5316 10140 5322 10192
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 6273 10115 6331 10121
rect 6273 10112 6285 10115
rect 5684 10084 6285 10112
rect 5684 10072 5690 10084
rect 6273 10081 6285 10084
rect 6319 10081 6331 10115
rect 6273 10075 6331 10081
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10044 5871 10047
rect 6086 10044 6092 10056
rect 5859 10016 6092 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 8312 10053 8340 10220
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 8757 10251 8815 10257
rect 8757 10217 8769 10251
rect 8803 10248 8815 10251
rect 9030 10248 9036 10260
rect 8803 10220 9036 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9398 10208 9404 10260
rect 9456 10208 9462 10260
rect 9674 10208 9680 10260
rect 9732 10208 9738 10260
rect 9766 10208 9772 10260
rect 9824 10208 9830 10260
rect 10686 10208 10692 10260
rect 10744 10208 10750 10260
rect 11238 10208 11244 10260
rect 11296 10208 11302 10260
rect 14645 10251 14703 10257
rect 14645 10217 14657 10251
rect 14691 10248 14703 10251
rect 18046 10248 18052 10260
rect 14691 10220 18052 10248
rect 14691 10217 14703 10220
rect 14645 10211 14703 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 20809 10251 20867 10257
rect 20809 10217 20821 10251
rect 20855 10248 20867 10251
rect 20898 10248 20904 10260
rect 20855 10220 20904 10248
rect 20855 10217 20867 10220
rect 20809 10211 20867 10217
rect 20898 10208 20904 10220
rect 20956 10208 20962 10260
rect 8386 10072 8392 10124
rect 8444 10072 8450 10124
rect 8570 10072 8576 10124
rect 8628 10112 8634 10124
rect 9033 10115 9091 10121
rect 9033 10112 9045 10115
rect 8628 10084 9045 10112
rect 8628 10072 8634 10084
rect 9033 10081 9045 10084
rect 9079 10081 9091 10115
rect 9033 10075 9091 10081
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10044 6239 10047
rect 8297 10047 8355 10053
rect 6227 10016 6316 10044
rect 6227 10013 6239 10016
rect 6181 10007 6239 10013
rect 6288 9988 6316 10016
rect 8297 10013 8309 10047
rect 8343 10013 8355 10047
rect 8297 10007 8355 10013
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9692 10044 9720 10208
rect 9171 10016 9720 10044
rect 9784 10044 9812 10208
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10112 10287 10115
rect 10502 10112 10508 10124
rect 10275 10084 10508 10112
rect 10275 10081 10287 10084
rect 10229 10075 10287 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10704 10112 10732 10208
rect 10965 10115 11023 10121
rect 10965 10112 10977 10115
rect 10704 10084 10977 10112
rect 10965 10081 10977 10084
rect 11011 10081 11023 10115
rect 10965 10075 11023 10081
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10112 11207 10115
rect 11256 10112 11284 10208
rect 19368 10183 19426 10189
rect 19368 10149 19380 10183
rect 19414 10180 19426 10183
rect 19797 10183 19855 10189
rect 19797 10180 19809 10183
rect 19414 10152 19809 10180
rect 19414 10149 19426 10152
rect 19368 10143 19426 10149
rect 19797 10149 19809 10152
rect 19843 10149 19855 10183
rect 19797 10143 19855 10149
rect 22738 10140 22744 10192
rect 22796 10140 22802 10192
rect 11195 10084 11284 10112
rect 11195 10081 11207 10084
rect 11149 10075 11207 10081
rect 14090 10072 14096 10124
rect 14148 10112 14154 10124
rect 14185 10115 14243 10121
rect 14185 10112 14197 10115
rect 14148 10084 14197 10112
rect 14148 10072 14154 10084
rect 14185 10081 14197 10084
rect 14231 10081 14243 10115
rect 14185 10075 14243 10081
rect 14458 10072 14464 10124
rect 14516 10072 14522 10124
rect 19610 10072 19616 10124
rect 19668 10072 19674 10124
rect 19702 10072 19708 10124
rect 19760 10072 19766 10124
rect 19886 10072 19892 10124
rect 19944 10072 19950 10124
rect 21085 10115 21143 10121
rect 21085 10081 21097 10115
rect 21131 10112 21143 10115
rect 21358 10112 21364 10124
rect 21131 10084 21364 10112
rect 21131 10081 21143 10084
rect 21085 10075 21143 10081
rect 21358 10072 21364 10084
rect 21416 10072 21422 10124
rect 21542 10072 21548 10124
rect 21600 10072 21606 10124
rect 21726 10072 21732 10124
rect 21784 10072 21790 10124
rect 22097 10115 22155 10121
rect 22097 10081 22109 10115
rect 22143 10112 22155 10115
rect 22756 10112 22784 10140
rect 22143 10084 22784 10112
rect 22143 10081 22155 10084
rect 22097 10075 22155 10081
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 9784 10016 10149 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 14274 10004 14280 10056
rect 14332 10004 14338 10056
rect 5626 9936 5632 9988
rect 5684 9936 5690 9988
rect 6270 9936 6276 9988
rect 6328 9936 6334 9988
rect 9490 9936 9496 9988
rect 9548 9976 9554 9988
rect 11698 9976 11704 9988
rect 9548 9948 11704 9976
rect 9548 9936 9554 9948
rect 11698 9936 11704 9948
rect 11756 9936 11762 9988
rect 4246 9868 4252 9920
rect 4304 9908 4310 9920
rect 5077 9911 5135 9917
rect 5077 9908 5089 9911
rect 4304 9880 5089 9908
rect 4304 9868 4310 9880
rect 5077 9877 5089 9880
rect 5123 9877 5135 9911
rect 5077 9871 5135 9877
rect 5261 9911 5319 9917
rect 5261 9877 5273 9911
rect 5307 9908 5319 9911
rect 6546 9908 6552 9920
rect 5307 9880 6552 9908
rect 5307 9877 5319 9880
rect 5261 9871 5319 9877
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 10594 9868 10600 9920
rect 10652 9868 10658 9920
rect 11146 9868 11152 9920
rect 11204 9868 11210 9920
rect 14182 9868 14188 9920
rect 14240 9868 14246 9920
rect 18233 9911 18291 9917
rect 18233 9877 18245 9911
rect 18279 9908 18291 9911
rect 18874 9908 18880 9920
rect 18279 9880 18880 9908
rect 18279 9877 18291 9880
rect 18233 9871 18291 9877
rect 18874 9868 18880 9880
rect 18932 9908 18938 9920
rect 19242 9908 19248 9920
rect 18932 9880 19248 9908
rect 18932 9868 18938 9880
rect 19242 9868 19248 9880
rect 19300 9868 19306 9920
rect 19720 9908 19748 10072
rect 20809 10047 20867 10053
rect 20809 10013 20821 10047
rect 20855 10044 20867 10047
rect 20898 10044 20904 10056
rect 20855 10016 20904 10044
rect 20855 10013 20867 10016
rect 20809 10007 20867 10013
rect 20898 10004 20904 10016
rect 20956 10044 20962 10056
rect 21821 10047 21879 10053
rect 21821 10044 21833 10047
rect 20956 10016 21833 10044
rect 20956 10004 20962 10016
rect 21821 10013 21833 10016
rect 21867 10013 21879 10047
rect 21821 10007 21879 10013
rect 20530 9936 20536 9988
rect 20588 9976 20594 9988
rect 21913 9979 21971 9985
rect 21913 9976 21925 9979
rect 20588 9948 21925 9976
rect 20588 9936 20594 9948
rect 21913 9945 21925 9948
rect 21959 9945 21971 9979
rect 21913 9939 21971 9945
rect 20622 9908 20628 9920
rect 19720 9880 20628 9908
rect 20622 9868 20628 9880
rect 20680 9908 20686 9920
rect 20993 9911 21051 9917
rect 20993 9908 21005 9911
rect 20680 9880 21005 9908
rect 20680 9868 20686 9880
rect 20993 9877 21005 9880
rect 21039 9877 21051 9911
rect 20993 9871 21051 9877
rect 21358 9868 21364 9920
rect 21416 9908 21422 9920
rect 22005 9911 22063 9917
rect 22005 9908 22017 9911
rect 21416 9880 22017 9908
rect 21416 9868 21422 9880
rect 22005 9877 22017 9880
rect 22051 9877 22063 9911
rect 22005 9871 22063 9877
rect 552 9818 23368 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 23368 9818
rect 552 9744 23368 9766
rect 5718 9664 5724 9716
rect 5776 9664 5782 9716
rect 6546 9664 6552 9716
rect 6604 9664 6610 9716
rect 7285 9707 7343 9713
rect 7285 9704 7297 9707
rect 7208 9676 7297 9704
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 7101 9639 7159 9645
rect 7101 9636 7113 9639
rect 5684 9608 7113 9636
rect 5684 9596 5690 9608
rect 7101 9605 7113 9608
rect 7147 9605 7159 9639
rect 7101 9599 7159 9605
rect 7208 9568 7236 9676
rect 7285 9673 7297 9676
rect 7331 9673 7343 9707
rect 7285 9667 7343 9673
rect 10594 9664 10600 9716
rect 10652 9704 10658 9716
rect 12069 9707 12127 9713
rect 12069 9704 12081 9707
rect 10652 9676 12081 9704
rect 10652 9664 10658 9676
rect 12069 9673 12081 9676
rect 12115 9673 12127 9707
rect 12069 9667 12127 9673
rect 14093 9707 14151 9713
rect 14093 9673 14105 9707
rect 14139 9704 14151 9707
rect 14182 9704 14188 9716
rect 14139 9676 14188 9704
rect 14139 9673 14151 9676
rect 14093 9667 14151 9673
rect 14182 9664 14188 9676
rect 14240 9664 14246 9716
rect 14274 9664 14280 9716
rect 14332 9664 14338 9716
rect 14458 9664 14464 9716
rect 14516 9664 14522 9716
rect 18325 9707 18383 9713
rect 18325 9673 18337 9707
rect 18371 9704 18383 9707
rect 19337 9707 19395 9713
rect 18371 9676 18460 9704
rect 18371 9673 18383 9676
rect 18325 9667 18383 9673
rect 11977 9639 12035 9645
rect 11977 9605 11989 9639
rect 12023 9636 12035 9639
rect 12529 9639 12587 9645
rect 12023 9608 12204 9636
rect 12023 9605 12035 9608
rect 11977 9599 12035 9605
rect 6012 9540 7236 9568
rect 10873 9571 10931 9577
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9500 4123 9503
rect 4246 9500 4252 9512
rect 4111 9472 4252 9500
rect 4111 9469 4123 9472
rect 4065 9463 4123 9469
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 4338 9460 4344 9512
rect 4396 9460 4402 9512
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 6012 9509 6040 9540
rect 5997 9503 6055 9509
rect 5997 9500 6009 9503
rect 5776 9472 6009 9500
rect 5776 9460 5782 9472
rect 5997 9469 6009 9472
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 6089 9503 6147 9509
rect 6089 9469 6101 9503
rect 6135 9500 6147 9503
rect 6178 9500 6184 9512
rect 6135 9472 6184 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 6748 9509 6776 9540
rect 10873 9537 10885 9571
rect 10919 9568 10931 9571
rect 11054 9568 11060 9580
rect 10919 9540 11060 9568
rect 10919 9537 10931 9540
rect 10873 9531 10931 9537
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 11146 9528 11152 9580
rect 11204 9568 11210 9580
rect 12176 9577 12204 9608
rect 12529 9605 12541 9639
rect 12575 9636 12587 9639
rect 14476 9636 14504 9664
rect 12575 9608 14504 9636
rect 18049 9639 18107 9645
rect 12575 9605 12587 9608
rect 12529 9599 12587 9605
rect 18049 9605 18061 9639
rect 18095 9636 18107 9639
rect 18230 9636 18236 9648
rect 18095 9608 18236 9636
rect 18095 9605 18107 9608
rect 18049 9599 18107 9605
rect 18230 9596 18236 9608
rect 18288 9596 18294 9648
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11204 9540 11529 9568
rect 11204 9528 11210 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 13633 9571 13691 9577
rect 13633 9568 13645 9571
rect 12860 9540 13645 9568
rect 12860 9528 12866 9540
rect 13633 9537 13645 9540
rect 13679 9537 13691 9571
rect 13633 9531 13691 9537
rect 14645 9571 14703 9577
rect 14645 9537 14657 9571
rect 14691 9568 14703 9571
rect 14826 9568 14832 9580
rect 14691 9540 14832 9568
rect 14691 9537 14703 9540
rect 14645 9531 14703 9537
rect 14826 9528 14832 9540
rect 14884 9528 14890 9580
rect 18432 9568 18460 9676
rect 19337 9673 19349 9707
rect 19383 9704 19395 9707
rect 19702 9704 19708 9716
rect 19383 9676 19708 9704
rect 19383 9673 19395 9676
rect 19337 9667 19395 9673
rect 19702 9664 19708 9676
rect 19760 9664 19766 9716
rect 19886 9664 19892 9716
rect 19944 9704 19950 9716
rect 20165 9707 20223 9713
rect 20165 9704 20177 9707
rect 19944 9676 20177 9704
rect 19944 9664 19950 9676
rect 20165 9673 20177 9676
rect 20211 9673 20223 9707
rect 20165 9667 20223 9673
rect 20714 9664 20720 9716
rect 20772 9664 20778 9716
rect 20806 9664 20812 9716
rect 20864 9704 20870 9716
rect 21085 9707 21143 9713
rect 21085 9704 21097 9707
rect 20864 9676 21097 9704
rect 20864 9664 20870 9676
rect 21085 9673 21097 9676
rect 21131 9704 21143 9707
rect 21726 9704 21732 9716
rect 21131 9676 21732 9704
rect 21131 9673 21143 9676
rect 21085 9667 21143 9673
rect 21726 9664 21732 9676
rect 21784 9664 21790 9716
rect 18509 9639 18567 9645
rect 18509 9605 18521 9639
rect 18555 9636 18567 9639
rect 20070 9636 20076 9648
rect 18555 9608 20076 9636
rect 18555 9605 18567 9608
rect 18509 9599 18567 9605
rect 20070 9596 20076 9608
rect 20128 9596 20134 9648
rect 20441 9639 20499 9645
rect 20441 9605 20453 9639
rect 20487 9605 20499 9639
rect 20441 9599 20499 9605
rect 20533 9639 20591 9645
rect 20533 9605 20545 9639
rect 20579 9636 20591 9639
rect 20732 9636 20760 9664
rect 20579 9608 20760 9636
rect 20579 9605 20591 9608
rect 20533 9599 20591 9605
rect 19242 9568 19248 9580
rect 18432 9540 19012 9568
rect 6733 9503 6791 9509
rect 6733 9469 6745 9503
rect 6779 9469 6791 9503
rect 6733 9463 6791 9469
rect 7006 9460 7012 9512
rect 7064 9460 7070 9512
rect 10962 9460 10968 9512
rect 11020 9460 11026 9512
rect 11609 9503 11667 9509
rect 11609 9469 11621 9503
rect 11655 9469 11667 9503
rect 11609 9463 11667 9469
rect 4586 9435 4644 9441
rect 4586 9432 4598 9435
rect 4264 9404 4598 9432
rect 4264 9373 4292 9404
rect 4586 9401 4598 9404
rect 4632 9401 4644 9435
rect 5813 9435 5871 9441
rect 5813 9432 5825 9435
rect 4586 9395 4644 9401
rect 5552 9404 5825 9432
rect 5552 9376 5580 9404
rect 5813 9401 5825 9404
rect 5859 9432 5871 9435
rect 6270 9432 6276 9444
rect 5859 9404 6276 9432
rect 5859 9401 5871 9404
rect 5813 9395 5871 9401
rect 6270 9392 6276 9404
rect 6328 9432 6334 9444
rect 6917 9435 6975 9441
rect 6917 9432 6929 9435
rect 6328 9404 6929 9432
rect 6328 9392 6334 9404
rect 6917 9401 6929 9404
rect 6963 9432 6975 9435
rect 7469 9435 7527 9441
rect 7469 9432 7481 9435
rect 6963 9404 7481 9432
rect 6963 9401 6975 9404
rect 6917 9395 6975 9401
rect 7469 9401 7481 9404
rect 7515 9401 7527 9435
rect 7469 9395 7527 9401
rect 11054 9392 11060 9444
rect 11112 9432 11118 9444
rect 11624 9432 11652 9463
rect 11698 9460 11704 9512
rect 11756 9500 11762 9512
rect 12345 9503 12403 9509
rect 12345 9500 12357 9503
rect 11756 9472 12357 9500
rect 11756 9460 11762 9472
rect 12345 9469 12357 9472
rect 12391 9469 12403 9503
rect 12345 9463 12403 9469
rect 13722 9460 13728 9512
rect 13780 9460 13786 9512
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 14240 9472 14565 9500
rect 14240 9460 14246 9472
rect 14553 9469 14565 9472
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 16393 9503 16451 9509
rect 16393 9469 16405 9503
rect 16439 9469 16451 9503
rect 16393 9463 16451 9469
rect 16577 9503 16635 9509
rect 16577 9469 16589 9503
rect 16623 9500 16635 9503
rect 16850 9500 16856 9512
rect 16623 9472 16856 9500
rect 16623 9469 16635 9472
rect 16577 9463 16635 9469
rect 11112 9404 11652 9432
rect 12069 9435 12127 9441
rect 11112 9392 11118 9404
rect 12069 9401 12081 9435
rect 12115 9401 12127 9435
rect 16408 9432 16436 9463
rect 16850 9460 16856 9472
rect 16908 9500 16914 9512
rect 17865 9503 17923 9509
rect 16908 9472 17816 9500
rect 16908 9460 16914 9472
rect 17678 9432 17684 9444
rect 16408 9404 17684 9432
rect 12069 9395 12127 9401
rect 4249 9367 4307 9373
rect 4249 9333 4261 9367
rect 4295 9333 4307 9367
rect 4249 9327 4307 9333
rect 5534 9324 5540 9376
rect 5592 9324 5598 9376
rect 5718 9324 5724 9376
rect 5776 9364 5782 9376
rect 6086 9364 6092 9376
rect 5776 9336 6092 9364
rect 5776 9324 5782 9336
rect 6086 9324 6092 9336
rect 6144 9364 6150 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 6144 9336 6193 9364
rect 6144 9324 6150 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6181 9327 6239 9333
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 6454 9364 6460 9376
rect 6411 9336 6460 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7259 9367 7317 9373
rect 7259 9364 7271 9367
rect 7064 9336 7271 9364
rect 7064 9324 7070 9336
rect 7259 9333 7271 9336
rect 7305 9333 7317 9367
rect 7259 9327 7317 9333
rect 11333 9367 11391 9373
rect 11333 9333 11345 9367
rect 11379 9364 11391 9367
rect 12084 9364 12112 9395
rect 17678 9392 17684 9404
rect 17736 9392 17742 9444
rect 17788 9432 17816 9472
rect 17865 9469 17877 9503
rect 17911 9500 17923 9503
rect 18690 9500 18696 9512
rect 17911 9472 18696 9500
rect 17911 9469 17923 9472
rect 17865 9463 17923 9469
rect 18690 9460 18696 9472
rect 18748 9460 18754 9512
rect 18782 9460 18788 9512
rect 18840 9460 18846 9512
rect 17788 9404 18092 9432
rect 11379 9336 12112 9364
rect 11379 9333 11391 9336
rect 11333 9327 11391 9333
rect 16482 9324 16488 9376
rect 16540 9324 16546 9376
rect 18064 9364 18092 9404
rect 18138 9392 18144 9444
rect 18196 9432 18202 9444
rect 18800 9432 18828 9460
rect 18984 9441 19012 9540
rect 19076 9540 19248 9568
rect 19076 9509 19104 9540
rect 19242 9528 19248 9540
rect 19300 9568 19306 9580
rect 20257 9571 20315 9577
rect 19300 9540 20024 9568
rect 19300 9528 19306 9540
rect 19061 9503 19119 9509
rect 19061 9469 19073 9503
rect 19107 9469 19119 9503
rect 19061 9463 19119 9469
rect 19334 9460 19340 9512
rect 19392 9460 19398 9512
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9469 19487 9503
rect 19429 9463 19487 9469
rect 18196 9404 18828 9432
rect 18969 9435 19027 9441
rect 18196 9392 18202 9404
rect 18969 9401 18981 9435
rect 19015 9432 19027 9435
rect 19352 9432 19380 9460
rect 19015 9404 19380 9432
rect 19444 9432 19472 9463
rect 19518 9460 19524 9512
rect 19576 9500 19582 9512
rect 19996 9509 20024 9540
rect 20257 9537 20269 9571
rect 20303 9568 20315 9571
rect 20349 9571 20407 9577
rect 20349 9568 20361 9571
rect 20303 9540 20361 9568
rect 20303 9537 20315 9540
rect 20257 9531 20315 9537
rect 20349 9537 20361 9540
rect 20395 9537 20407 9571
rect 20456 9568 20484 9599
rect 22554 9596 22560 9648
rect 22612 9596 22618 9648
rect 22465 9571 22523 9577
rect 20456 9540 21220 9568
rect 20349 9531 20407 9537
rect 19705 9503 19763 9509
rect 19705 9500 19717 9503
rect 19576 9472 19717 9500
rect 19576 9460 19582 9472
rect 19705 9469 19717 9472
rect 19751 9469 19763 9503
rect 19705 9463 19763 9469
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9469 20039 9503
rect 19981 9463 20039 9469
rect 20162 9460 20168 9512
rect 20220 9500 20226 9512
rect 20272 9500 20300 9531
rect 20220 9472 20484 9500
rect 20220 9460 20226 9472
rect 20346 9432 20352 9444
rect 19444 9404 20352 9432
rect 19015 9401 19027 9404
rect 18969 9395 19027 9401
rect 18341 9367 18399 9373
rect 18341 9364 18353 9367
rect 18064 9336 18353 9364
rect 18341 9333 18353 9336
rect 18387 9364 18399 9367
rect 19153 9367 19211 9373
rect 19153 9364 19165 9367
rect 18387 9336 19165 9364
rect 18387 9333 18399 9336
rect 18341 9327 18399 9333
rect 19153 9333 19165 9336
rect 19199 9364 19211 9367
rect 19444 9364 19472 9404
rect 20346 9392 20352 9404
rect 20404 9392 20410 9444
rect 19199 9336 19472 9364
rect 19521 9367 19579 9373
rect 19199 9333 19211 9336
rect 19153 9327 19211 9333
rect 19521 9333 19533 9367
rect 19567 9364 19579 9367
rect 19702 9364 19708 9376
rect 19567 9336 19708 9364
rect 19567 9333 19579 9336
rect 19521 9327 19579 9333
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 19889 9367 19947 9373
rect 19889 9333 19901 9367
rect 19935 9364 19947 9367
rect 20162 9364 20168 9376
rect 19935 9336 20168 9364
rect 19935 9333 19947 9336
rect 19889 9327 19947 9333
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 20456 9364 20484 9472
rect 20622 9460 20628 9512
rect 20680 9460 20686 9512
rect 20717 9503 20775 9509
rect 20717 9469 20729 9503
rect 20763 9500 20775 9503
rect 21082 9500 21088 9512
rect 20763 9472 21088 9500
rect 20763 9469 20775 9472
rect 20717 9463 20775 9469
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 21192 9500 21220 9540
rect 22465 9537 22477 9571
rect 22511 9568 22523 9571
rect 22572 9568 22600 9596
rect 22511 9540 22600 9568
rect 22511 9537 22523 9540
rect 22465 9531 22523 9537
rect 22557 9503 22615 9509
rect 22557 9500 22569 9503
rect 21192 9472 22569 9500
rect 22557 9469 22569 9472
rect 22603 9469 22615 9503
rect 22557 9463 22615 9469
rect 22741 9503 22799 9509
rect 22741 9469 22753 9503
rect 22787 9469 22799 9503
rect 22741 9463 22799 9469
rect 21358 9432 21364 9444
rect 20824 9404 21364 9432
rect 20824 9376 20852 9404
rect 21358 9392 21364 9404
rect 21416 9392 21422 9444
rect 22220 9435 22278 9441
rect 22220 9401 22232 9435
rect 22266 9432 22278 9435
rect 22649 9435 22707 9441
rect 22649 9432 22661 9435
rect 22266 9404 22661 9432
rect 22266 9401 22278 9404
rect 22220 9395 22278 9401
rect 22649 9401 22661 9404
rect 22695 9401 22707 9435
rect 22649 9395 22707 9401
rect 20714 9364 20720 9376
rect 20456 9336 20720 9364
rect 20714 9324 20720 9336
rect 20772 9324 20778 9376
rect 20806 9324 20812 9376
rect 20864 9324 20870 9376
rect 20898 9324 20904 9376
rect 20956 9324 20962 9376
rect 21376 9364 21404 9392
rect 22094 9364 22100 9376
rect 21376 9336 22100 9364
rect 22094 9324 22100 9336
rect 22152 9364 22158 9376
rect 22756 9364 22784 9463
rect 22152 9336 22784 9364
rect 22152 9324 22158 9336
rect 552 9274 23368 9296
rect 552 9222 19022 9274
rect 19074 9222 19086 9274
rect 19138 9222 19150 9274
rect 19202 9222 19214 9274
rect 19266 9222 19278 9274
rect 19330 9222 23368 9274
rect 552 9200 23368 9222
rect 4338 9120 4344 9172
rect 4396 9120 4402 9172
rect 5813 9163 5871 9169
rect 5813 9129 5825 9163
rect 5859 9160 5871 9163
rect 6178 9160 6184 9172
rect 5859 9132 6184 9160
rect 5859 9129 5871 9132
rect 5813 9123 5871 9129
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 6454 9120 6460 9172
rect 6512 9160 6518 9172
rect 8037 9163 8095 9169
rect 8037 9160 8049 9163
rect 6512 9132 8049 9160
rect 6512 9120 6518 9132
rect 8037 9129 8049 9132
rect 8083 9160 8095 9163
rect 8754 9160 8760 9172
rect 8083 9132 8760 9160
rect 8083 9129 8095 9132
rect 8037 9123 8095 9129
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 14090 9120 14096 9172
rect 14148 9160 14154 9172
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 14148 9132 14197 9160
rect 14148 9120 14154 9132
rect 14185 9129 14197 9132
rect 14231 9129 14243 9163
rect 14185 9123 14243 9129
rect 16482 9120 16488 9172
rect 16540 9120 16546 9172
rect 17310 9120 17316 9172
rect 17368 9160 17374 9172
rect 17497 9163 17555 9169
rect 17497 9160 17509 9163
rect 17368 9132 17509 9160
rect 17368 9120 17374 9132
rect 17497 9129 17509 9132
rect 17543 9129 17555 9163
rect 17497 9123 17555 9129
rect 17865 9163 17923 9169
rect 17865 9129 17877 9163
rect 17911 9160 17923 9163
rect 17954 9160 17960 9172
rect 17911 9132 17960 9160
rect 17911 9129 17923 9132
rect 17865 9123 17923 9129
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 18230 9120 18236 9172
rect 18288 9120 18294 9172
rect 18690 9120 18696 9172
rect 18748 9160 18754 9172
rect 19613 9163 19671 9169
rect 19613 9160 19625 9163
rect 18748 9132 19625 9160
rect 18748 9120 18754 9132
rect 19613 9129 19625 9132
rect 19659 9129 19671 9163
rect 20717 9163 20775 9169
rect 20717 9160 20729 9163
rect 19613 9123 19671 9129
rect 19812 9132 20729 9160
rect 4356 9092 4384 9120
rect 7098 9092 7104 9104
rect 4356 9064 7104 9092
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 4356 9024 4384 9064
rect 7098 9052 7104 9064
rect 7156 9092 7162 9104
rect 7156 9064 7236 9092
rect 7156 9052 7162 9064
rect 4295 8996 4384 9024
rect 4516 9027 4574 9033
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 4516 8993 4528 9027
rect 4562 9024 4574 9027
rect 4890 9024 4896 9036
rect 4562 8996 4896 9024
rect 4562 8993 4574 8996
rect 4516 8987 4574 8993
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 6362 8984 6368 9036
rect 6420 9024 6426 9036
rect 7208 9033 7236 9064
rect 7742 9052 7748 9104
rect 7800 9092 7806 9104
rect 7837 9095 7895 9101
rect 7837 9092 7849 9095
rect 7800 9064 7849 9092
rect 7800 9052 7806 9064
rect 7837 9061 7849 9064
rect 7883 9061 7895 9095
rect 14918 9092 14924 9104
rect 7837 9055 7895 9061
rect 13832 9064 14924 9092
rect 13832 9033 13860 9064
rect 14918 9052 14924 9064
rect 14976 9052 14982 9104
rect 16384 9095 16442 9101
rect 16384 9061 16396 9095
rect 16430 9092 16442 9095
rect 16500 9092 16528 9120
rect 16430 9064 16528 9092
rect 18248 9092 18276 9120
rect 19812 9104 19840 9132
rect 20717 9129 20729 9132
rect 20763 9129 20775 9163
rect 20898 9160 20904 9172
rect 20717 9123 20775 9129
rect 20824 9132 20904 9160
rect 18386 9095 18444 9101
rect 18386 9092 18398 9095
rect 18248 9064 18398 9092
rect 16430 9061 16442 9064
rect 16384 9055 16442 9061
rect 18386 9061 18398 9064
rect 18432 9061 18444 9095
rect 18386 9055 18444 9061
rect 18782 9052 18788 9104
rect 18840 9092 18846 9104
rect 19702 9092 19708 9104
rect 18840 9064 19708 9092
rect 18840 9052 18846 9064
rect 19702 9052 19708 9064
rect 19760 9052 19766 9104
rect 19794 9052 19800 9104
rect 19852 9052 19858 9104
rect 20533 9095 20591 9101
rect 20533 9092 20545 9095
rect 19996 9064 20545 9092
rect 6926 9027 6984 9033
rect 6926 9024 6938 9027
rect 6420 8996 6938 9024
rect 6420 8984 6426 8996
rect 6926 8993 6938 8996
rect 6972 8993 6984 9027
rect 6926 8987 6984 8993
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 8993 7251 9027
rect 7193 8987 7251 8993
rect 13173 9027 13231 9033
rect 13173 8993 13185 9027
rect 13219 8993 13231 9027
rect 13173 8987 13231 8993
rect 13817 9027 13875 9033
rect 13817 8993 13829 9027
rect 13863 8993 13875 9027
rect 13817 8987 13875 8993
rect 13188 8888 13216 8987
rect 16850 8984 16856 9036
rect 16908 9024 16914 9036
rect 17773 9027 17831 9033
rect 17773 9024 17785 9027
rect 16908 8996 17785 9024
rect 16908 8984 16914 8996
rect 17773 8993 17785 8996
rect 17819 8993 17831 9027
rect 17773 8987 17831 8993
rect 18049 9027 18107 9033
rect 18049 8993 18061 9027
rect 18095 9024 18107 9027
rect 19996 9024 20024 9064
rect 20533 9061 20545 9064
rect 20579 9061 20591 9095
rect 20533 9055 20591 9061
rect 18095 8996 20024 9024
rect 18095 8993 18107 8996
rect 18049 8987 18107 8993
rect 20070 8984 20076 9036
rect 20128 9024 20134 9036
rect 20165 9027 20223 9033
rect 20165 9024 20177 9027
rect 20128 8996 20177 9024
rect 20128 8984 20134 8996
rect 20165 8993 20177 8996
rect 20211 8993 20223 9027
rect 20165 8987 20223 8993
rect 20257 9027 20315 9033
rect 20257 8993 20269 9027
rect 20303 8993 20315 9027
rect 20257 8987 20315 8993
rect 13906 8916 13912 8968
rect 13964 8916 13970 8968
rect 16117 8959 16175 8965
rect 16117 8925 16129 8959
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 14550 8888 14556 8900
rect 8036 8860 8616 8888
rect 13188 8860 14556 8888
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 5534 8820 5540 8832
rect 5224 8792 5540 8820
rect 5224 8780 5230 8792
rect 5534 8780 5540 8792
rect 5592 8820 5598 8832
rect 5629 8823 5687 8829
rect 5629 8820 5641 8823
rect 5592 8792 5641 8820
rect 5592 8780 5598 8792
rect 5629 8789 5641 8792
rect 5675 8789 5687 8823
rect 5629 8783 5687 8789
rect 5810 8780 5816 8832
rect 5868 8820 5874 8832
rect 7558 8820 7564 8832
rect 5868 8792 7564 8820
rect 5868 8780 5874 8792
rect 7558 8780 7564 8792
rect 7616 8820 7622 8832
rect 7926 8820 7932 8832
rect 7616 8792 7932 8820
rect 7616 8780 7622 8792
rect 7926 8780 7932 8792
rect 7984 8780 7990 8832
rect 8036 8829 8064 8860
rect 8588 8832 8616 8860
rect 14550 8848 14556 8860
rect 14608 8848 14614 8900
rect 16132 8832 16160 8919
rect 18138 8916 18144 8968
rect 18196 8916 18202 8968
rect 19426 8916 19432 8968
rect 19484 8916 19490 8968
rect 19518 8916 19524 8968
rect 19576 8916 19582 8968
rect 19702 8916 19708 8968
rect 19760 8956 19766 8968
rect 20272 8956 20300 8987
rect 20346 8984 20352 9036
rect 20404 8984 20410 9036
rect 20824 9024 20852 9132
rect 20898 9120 20904 9132
rect 20956 9120 20962 9172
rect 21082 9120 21088 9172
rect 21140 9120 21146 9172
rect 21266 9120 21272 9172
rect 21324 9160 21330 9172
rect 22554 9160 22560 9172
rect 21324 9132 22560 9160
rect 21324 9120 21330 9132
rect 22554 9120 22560 9132
rect 22612 9120 22618 9172
rect 22649 9163 22707 9169
rect 22649 9129 22661 9163
rect 22695 9160 22707 9163
rect 22738 9160 22744 9172
rect 22695 9132 22744 9160
rect 22695 9129 22707 9132
rect 22649 9123 22707 9129
rect 22738 9120 22744 9132
rect 22796 9120 22802 9172
rect 21100 9092 21128 9120
rect 20916 9064 22784 9092
rect 20916 9033 20944 9064
rect 20548 8996 20852 9024
rect 20901 9027 20959 9033
rect 20548 8965 20576 8996
rect 20901 8993 20913 9027
rect 20947 8993 20959 9027
rect 21525 9027 21583 9033
rect 21525 9024 21537 9027
rect 20901 8987 20959 8993
rect 21100 8996 21537 9024
rect 19760 8928 20300 8956
rect 20533 8959 20591 8965
rect 19760 8916 19766 8928
rect 20533 8925 20545 8959
rect 20579 8925 20591 8959
rect 21100 8956 21128 8996
rect 21525 8993 21537 8996
rect 21571 8993 21583 9027
rect 21525 8987 21583 8993
rect 22002 8984 22008 9036
rect 22060 9024 22066 9036
rect 22756 9033 22784 9064
rect 22741 9027 22799 9033
rect 22060 8996 22508 9024
rect 22060 8984 22066 8996
rect 20533 8919 20591 8925
rect 20640 8928 21128 8956
rect 17052 8860 18184 8888
rect 8021 8823 8079 8829
rect 8021 8789 8033 8823
rect 8067 8789 8079 8823
rect 8021 8783 8079 8789
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 8205 8823 8263 8829
rect 8205 8820 8217 8823
rect 8168 8792 8217 8820
rect 8168 8780 8174 8792
rect 8205 8789 8217 8792
rect 8251 8789 8263 8823
rect 8205 8783 8263 8789
rect 8570 8780 8576 8832
rect 8628 8780 8634 8832
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 13357 8823 13415 8829
rect 13357 8820 13369 8823
rect 9640 8792 13369 8820
rect 9640 8780 9646 8792
rect 13357 8789 13369 8792
rect 13403 8820 13415 8823
rect 14458 8820 14464 8832
rect 13403 8792 14464 8820
rect 13403 8789 13415 8792
rect 13357 8783 13415 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 16114 8780 16120 8832
rect 16172 8820 16178 8832
rect 17052 8820 17080 8860
rect 16172 8792 17080 8820
rect 16172 8780 16178 8792
rect 18046 8780 18052 8832
rect 18104 8780 18110 8832
rect 18156 8820 18184 8860
rect 19444 8820 19472 8916
rect 19536 8829 19564 8916
rect 19978 8848 19984 8900
rect 20036 8888 20042 8900
rect 20548 8888 20576 8919
rect 20036 8860 20576 8888
rect 20036 8848 20042 8860
rect 20640 8832 20668 8928
rect 21266 8916 21272 8968
rect 21324 8916 21330 8968
rect 22480 8956 22508 8996
rect 22741 8993 22753 9027
rect 22787 8993 22799 9027
rect 22741 8987 22799 8993
rect 22480 8928 22968 8956
rect 22940 8897 22968 8928
rect 22925 8891 22983 8897
rect 22925 8857 22937 8891
rect 22971 8857 22983 8891
rect 22925 8851 22983 8857
rect 18156 8792 19472 8820
rect 19521 8823 19579 8829
rect 19521 8789 19533 8823
rect 19567 8789 19579 8823
rect 19521 8783 19579 8789
rect 19797 8823 19855 8829
rect 19797 8789 19809 8823
rect 19843 8820 19855 8823
rect 20162 8820 20168 8832
rect 19843 8792 20168 8820
rect 19843 8789 19855 8792
rect 19797 8783 19855 8789
rect 20162 8780 20168 8792
rect 20220 8780 20226 8832
rect 20622 8780 20628 8832
rect 20680 8780 20686 8832
rect 552 8730 23368 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 23368 8730
rect 552 8656 23368 8678
rect 4890 8576 4896 8628
rect 4948 8576 4954 8628
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5350 8616 5356 8628
rect 5132 8588 5356 8616
rect 5132 8576 5138 8588
rect 5350 8576 5356 8588
rect 5408 8616 5414 8628
rect 5408 8588 5580 8616
rect 5408 8576 5414 8588
rect 5445 8551 5503 8557
rect 5445 8548 5457 8551
rect 4908 8520 5457 8548
rect 4908 8421 4936 8520
rect 5445 8517 5457 8520
rect 5491 8517 5503 8551
rect 5552 8548 5580 8588
rect 5626 8576 5632 8628
rect 5684 8616 5690 8628
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5684 8588 6009 8616
rect 5684 8576 5690 8588
rect 5997 8585 6009 8588
rect 6043 8585 6055 8619
rect 5997 8579 6055 8585
rect 6178 8576 6184 8628
rect 6236 8576 6242 8628
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 6362 8616 6368 8628
rect 6319 8588 6368 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 7208 8588 7696 8616
rect 5718 8548 5724 8560
rect 5552 8520 5724 8548
rect 5445 8511 5503 8517
rect 5718 8508 5724 8520
rect 5776 8508 5782 8560
rect 5810 8508 5816 8560
rect 5868 8508 5874 8560
rect 6196 8548 6224 8576
rect 5920 8520 6224 8548
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 5828 8480 5856 8508
rect 5583 8452 5856 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 4893 8415 4951 8421
rect 4893 8381 4905 8415
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 5074 8372 5080 8424
rect 5132 8412 5138 8424
rect 5920 8421 5948 8520
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8480 6239 8483
rect 7208 8480 7236 8588
rect 7282 8508 7288 8560
rect 7340 8508 7346 8560
rect 7558 8548 7564 8560
rect 7484 8520 7564 8548
rect 6227 8452 7236 8480
rect 7377 8483 7435 8489
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 7377 8449 7389 8483
rect 7423 8480 7435 8483
rect 7484 8480 7512 8520
rect 7558 8508 7564 8520
rect 7616 8508 7622 8560
rect 7668 8548 7696 8588
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 10134 8616 10140 8628
rect 7984 8588 10140 8616
rect 7984 8576 7990 8588
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 14734 8616 14740 8628
rect 10244 8588 11560 8616
rect 8294 8548 8300 8560
rect 7668 8520 8300 8548
rect 8294 8508 8300 8520
rect 8352 8548 8358 8560
rect 10244 8548 10272 8588
rect 8352 8520 10272 8548
rect 8352 8508 8358 8520
rect 7423 8452 7512 8480
rect 7576 8452 7788 8480
rect 7423 8449 7435 8452
rect 7377 8443 7435 8449
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 5132 8384 5181 8412
rect 5132 8372 5138 8384
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 5905 8415 5963 8421
rect 5169 8375 5227 8381
rect 5271 8393 5329 8399
rect 5271 8359 5283 8393
rect 5317 8378 5329 8393
rect 5905 8381 5917 8415
rect 5951 8381 5963 8415
rect 5317 8359 5396 8378
rect 5905 8375 5963 8381
rect 6273 8415 6331 8421
rect 6273 8381 6285 8415
rect 6319 8381 6331 8415
rect 6273 8375 6331 8381
rect 5271 8353 5396 8359
rect 5276 8350 5396 8353
rect 5077 8279 5135 8285
rect 5077 8245 5089 8279
rect 5123 8276 5135 8279
rect 5166 8276 5172 8288
rect 5123 8248 5172 8276
rect 5123 8245 5135 8248
rect 5077 8239 5135 8245
rect 5166 8236 5172 8248
rect 5224 8276 5230 8288
rect 5368 8276 5396 8350
rect 6181 8347 6239 8353
rect 6181 8313 6193 8347
rect 6227 8344 6239 8347
rect 6288 8344 6316 8375
rect 6454 8372 6460 8424
rect 6512 8412 6518 8424
rect 7576 8421 7604 8452
rect 7760 8421 7788 8452
rect 8202 8440 8208 8492
rect 8260 8440 8266 8492
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8444 8452 8708 8480
rect 8444 8440 8450 8452
rect 7009 8415 7067 8421
rect 7009 8412 7021 8415
rect 6512 8384 7021 8412
rect 6512 8372 6518 8384
rect 7009 8381 7021 8384
rect 7055 8412 7067 8415
rect 7561 8415 7619 8421
rect 7561 8412 7573 8415
rect 7055 8384 7573 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 7561 8381 7573 8384
rect 7607 8381 7619 8415
rect 7561 8375 7619 8381
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8381 7711 8415
rect 7653 8375 7711 8381
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8381 7803 8415
rect 7745 8375 7803 8381
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8412 8079 8415
rect 8570 8412 8576 8424
rect 8067 8384 8576 8412
rect 8067 8381 8079 8384
rect 8021 8375 8079 8381
rect 6227 8316 6316 8344
rect 7285 8347 7343 8353
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 7285 8313 7297 8347
rect 7331 8344 7343 8347
rect 7377 8347 7435 8353
rect 7377 8344 7389 8347
rect 7331 8316 7389 8344
rect 7331 8313 7343 8316
rect 7285 8307 7343 8313
rect 7377 8313 7389 8316
rect 7423 8313 7435 8347
rect 7377 8307 7435 8313
rect 5224 8248 5396 8276
rect 7101 8279 7159 8285
rect 5224 8236 5230 8248
rect 7101 8245 7113 8279
rect 7147 8276 7159 8279
rect 7668 8276 7696 8375
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8680 8421 8708 8452
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 10134 8440 10140 8492
rect 10192 8480 10198 8492
rect 10229 8483 10287 8489
rect 10229 8480 10241 8483
rect 10192 8452 10241 8480
rect 10192 8440 10198 8452
rect 10229 8449 10241 8452
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 10778 8480 10784 8492
rect 10459 8452 10784 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8381 8723 8415
rect 8665 8375 8723 8381
rect 8772 8353 8800 8440
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8412 8999 8415
rect 9030 8412 9036 8424
rect 8987 8384 9036 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9030 8372 9036 8384
rect 9088 8412 9094 8424
rect 10428 8412 10456 8443
rect 10778 8440 10784 8452
rect 10836 8480 10842 8492
rect 11532 8489 11560 8588
rect 13924 8588 14740 8616
rect 12526 8508 12532 8560
rect 12584 8548 12590 8560
rect 13541 8551 13599 8557
rect 13541 8548 13553 8551
rect 12584 8520 13553 8548
rect 12584 8508 12590 8520
rect 13541 8517 13553 8520
rect 13587 8548 13599 8551
rect 13722 8548 13728 8560
rect 13587 8520 13728 8548
rect 13587 8517 13599 8520
rect 13541 8511 13599 8517
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 11517 8483 11575 8489
rect 10836 8452 11192 8480
rect 10836 8440 10842 8452
rect 9088 8384 10456 8412
rect 9088 8372 9094 8384
rect 10502 8372 10508 8424
rect 10560 8372 10566 8424
rect 10962 8372 10968 8424
rect 11020 8412 11026 8424
rect 11164 8421 11192 8452
rect 11517 8449 11529 8483
rect 11563 8480 11575 8483
rect 13630 8480 13636 8492
rect 11563 8452 13636 8480
rect 11563 8449 11575 8452
rect 11517 8443 11575 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 11057 8415 11115 8421
rect 11057 8412 11069 8415
rect 11020 8384 11069 8412
rect 11020 8372 11026 8384
rect 11057 8381 11069 8384
rect 11103 8381 11115 8415
rect 11057 8375 11115 8381
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 8389 8347 8447 8353
rect 8389 8344 8401 8347
rect 8312 8316 8401 8344
rect 7742 8276 7748 8288
rect 7147 8248 7748 8276
rect 7147 8245 7159 8248
rect 7101 8239 7159 8245
rect 7742 8236 7748 8248
rect 7800 8276 7806 8288
rect 7837 8279 7895 8285
rect 7837 8276 7849 8279
rect 7800 8248 7849 8276
rect 7800 8236 7806 8248
rect 7837 8245 7849 8248
rect 7883 8276 7895 8279
rect 8312 8276 8340 8316
rect 8389 8313 8401 8316
rect 8435 8313 8447 8347
rect 8389 8307 8447 8313
rect 8757 8347 8815 8353
rect 8757 8313 8769 8347
rect 8803 8313 8815 8347
rect 10520 8344 10548 8372
rect 10686 8344 10692 8356
rect 10520 8316 10692 8344
rect 8757 8307 8815 8313
rect 10686 8304 10692 8316
rect 10744 8344 10750 8356
rect 10781 8347 10839 8353
rect 10781 8344 10793 8347
rect 10744 8316 10793 8344
rect 10744 8304 10750 8316
rect 10781 8313 10793 8316
rect 10827 8313 10839 8347
rect 11072 8344 11100 8375
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 11296 8384 11713 8412
rect 11296 8372 11302 8384
rect 11701 8381 11713 8384
rect 11747 8381 11759 8415
rect 11701 8375 11759 8381
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8381 11851 8415
rect 11793 8375 11851 8381
rect 12529 8415 12587 8421
rect 12529 8381 12541 8415
rect 12575 8412 12587 8415
rect 13170 8412 13176 8424
rect 12575 8384 13176 8412
rect 12575 8381 12587 8384
rect 12529 8375 12587 8381
rect 11808 8344 11836 8375
rect 13170 8372 13176 8384
rect 13228 8372 13234 8424
rect 13924 8421 13952 8588
rect 14734 8576 14740 8588
rect 14792 8576 14798 8628
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 15841 8619 15899 8625
rect 15841 8616 15853 8619
rect 15611 8588 15853 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 15841 8585 15853 8588
rect 15887 8585 15899 8619
rect 15841 8579 15899 8585
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 17218 8616 17224 8628
rect 16724 8588 17224 8616
rect 16724 8576 16730 8588
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 17678 8576 17684 8628
rect 17736 8576 17742 8628
rect 18046 8576 18052 8628
rect 18104 8576 18110 8628
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 18690 8616 18696 8628
rect 18196 8588 18696 8616
rect 18196 8576 18202 8588
rect 18690 8576 18696 8588
rect 18748 8616 18754 8628
rect 19610 8616 19616 8628
rect 18748 8588 19616 8616
rect 18748 8576 18754 8588
rect 19610 8576 19616 8588
rect 19668 8576 19674 8628
rect 19702 8576 19708 8628
rect 19760 8616 19766 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 19760 8588 20085 8616
rect 19760 8576 19766 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 20073 8579 20131 8585
rect 20622 8576 20628 8628
rect 20680 8576 20686 8628
rect 21085 8619 21143 8625
rect 21085 8585 21097 8619
rect 21131 8616 21143 8619
rect 21361 8619 21419 8625
rect 21361 8616 21373 8619
rect 21131 8588 21373 8616
rect 21131 8585 21143 8588
rect 21085 8579 21143 8585
rect 21361 8585 21373 8588
rect 21407 8585 21419 8619
rect 21361 8579 21419 8585
rect 21818 8576 21824 8628
rect 21876 8616 21882 8628
rect 22189 8619 22247 8625
rect 22189 8616 22201 8619
rect 21876 8588 22201 8616
rect 21876 8576 21882 8588
rect 22189 8585 22201 8588
rect 22235 8585 22247 8619
rect 22189 8579 22247 8585
rect 13998 8508 14004 8560
rect 14056 8548 14062 8560
rect 14093 8551 14151 8557
rect 14093 8548 14105 8551
rect 14056 8520 14105 8548
rect 14056 8508 14062 8520
rect 14093 8517 14105 8520
rect 14139 8548 14151 8551
rect 14139 8520 15148 8548
rect 14139 8517 14151 8520
rect 14093 8511 14151 8517
rect 14642 8440 14648 8492
rect 14700 8440 14706 8492
rect 15120 8424 15148 8520
rect 15654 8508 15660 8560
rect 15712 8508 15718 8560
rect 16022 8508 16028 8560
rect 16080 8508 16086 8560
rect 16209 8551 16267 8557
rect 16209 8517 16221 8551
rect 16255 8548 16267 8551
rect 17037 8551 17095 8557
rect 17037 8548 17049 8551
rect 16255 8520 17049 8548
rect 16255 8517 16267 8520
rect 16209 8511 16267 8517
rect 17037 8517 17049 8520
rect 17083 8548 17095 8551
rect 17589 8551 17647 8557
rect 17589 8548 17601 8551
rect 17083 8520 17601 8548
rect 17083 8517 17095 8520
rect 17037 8511 17095 8517
rect 17589 8517 17601 8520
rect 17635 8517 17647 8551
rect 17862 8548 17868 8560
rect 17589 8511 17647 8517
rect 17788 8520 17868 8548
rect 16040 8480 16068 8508
rect 16301 8483 16359 8489
rect 16301 8480 16313 8483
rect 15212 8452 16313 8480
rect 13909 8415 13967 8421
rect 13909 8381 13921 8415
rect 13955 8381 13967 8415
rect 13909 8375 13967 8381
rect 14458 8372 14464 8424
rect 14516 8372 14522 8424
rect 14826 8372 14832 8424
rect 14884 8372 14890 8424
rect 14921 8415 14979 8421
rect 14921 8381 14933 8415
rect 14967 8381 14979 8415
rect 14921 8375 14979 8381
rect 11072 8316 11836 8344
rect 13817 8347 13875 8353
rect 10781 8307 10839 8313
rect 13817 8313 13829 8347
rect 13863 8344 13875 8347
rect 13863 8316 14504 8344
rect 13863 8313 13875 8316
rect 13817 8307 13875 8313
rect 7883 8248 8340 8276
rect 7883 8245 7895 8248
rect 7837 8239 7895 8245
rect 10226 8236 10232 8288
rect 10284 8236 10290 8288
rect 10502 8236 10508 8288
rect 10560 8276 10566 8288
rect 10965 8279 11023 8285
rect 10965 8276 10977 8279
rect 10560 8248 10977 8276
rect 10560 8236 10566 8248
rect 10965 8245 10977 8248
rect 11011 8276 11023 8279
rect 11054 8276 11060 8288
rect 11011 8248 11060 8276
rect 11011 8245 11023 8248
rect 10965 8239 11023 8245
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 11330 8236 11336 8288
rect 11388 8236 11394 8288
rect 11517 8279 11575 8285
rect 11517 8245 11529 8279
rect 11563 8276 11575 8279
rect 11606 8276 11612 8288
rect 11563 8248 11612 8276
rect 11563 8245 11575 8248
rect 11517 8239 11575 8245
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 12710 8236 12716 8288
rect 12768 8236 12774 8288
rect 13722 8236 13728 8288
rect 13780 8236 13786 8288
rect 14366 8236 14372 8288
rect 14424 8236 14430 8288
rect 14476 8276 14504 8316
rect 14642 8304 14648 8356
rect 14700 8304 14706 8356
rect 14936 8288 14964 8375
rect 15102 8372 15108 8424
rect 15160 8372 15166 8424
rect 15212 8421 15240 8452
rect 16301 8449 16313 8452
rect 16347 8449 16359 8483
rect 16666 8480 16672 8492
rect 16301 8443 16359 8449
rect 16500 8452 16672 8480
rect 16500 8421 16528 8452
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 16850 8440 16856 8492
rect 16908 8440 16914 8492
rect 17310 8440 17316 8492
rect 17368 8440 17374 8492
rect 17788 8489 17816 8520
rect 17862 8508 17868 8520
rect 17920 8508 17926 8560
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8449 17831 8483
rect 18064 8480 18092 8576
rect 20806 8548 20812 8560
rect 20364 8520 20812 8548
rect 18064 8452 18828 8480
rect 17773 8443 17831 8449
rect 15197 8415 15255 8421
rect 15197 8381 15209 8415
rect 15243 8381 15255 8415
rect 15197 8375 15255 8381
rect 15381 8415 15439 8421
rect 15381 8381 15393 8415
rect 15427 8412 15439 8415
rect 16485 8415 16543 8421
rect 16485 8412 16497 8415
rect 15427 8384 16497 8412
rect 15427 8381 15439 8384
rect 15381 8375 15439 8381
rect 16485 8381 16497 8384
rect 16531 8381 16543 8415
rect 16485 8375 16543 8381
rect 16577 8415 16635 8421
rect 16577 8381 16589 8415
rect 16623 8412 16635 8415
rect 17328 8412 17356 8440
rect 17497 8415 17555 8421
rect 17497 8412 17509 8415
rect 16623 8384 17509 8412
rect 16623 8381 16635 8384
rect 16577 8375 16635 8381
rect 17497 8381 17509 8384
rect 17543 8381 17555 8415
rect 17497 8375 17555 8381
rect 18690 8372 18696 8424
rect 18748 8372 18754 8424
rect 18800 8412 18828 8452
rect 20364 8421 20392 8520
rect 20806 8508 20812 8520
rect 20864 8508 20870 8560
rect 21269 8551 21327 8557
rect 21269 8517 21281 8551
rect 21315 8548 21327 8551
rect 21315 8520 22508 8548
rect 21315 8517 21327 8520
rect 21269 8511 21327 8517
rect 20456 8452 20852 8480
rect 20456 8421 20484 8452
rect 18949 8415 19007 8421
rect 18949 8412 18961 8415
rect 18800 8384 18961 8412
rect 18949 8381 18961 8384
rect 18995 8381 19007 8415
rect 18949 8375 19007 8381
rect 20349 8415 20407 8421
rect 20349 8381 20361 8415
rect 20395 8381 20407 8415
rect 20349 8375 20407 8381
rect 20441 8415 20499 8421
rect 20441 8381 20453 8415
rect 20487 8381 20499 8415
rect 20441 8375 20499 8381
rect 20530 8372 20536 8424
rect 20588 8412 20594 8424
rect 20625 8415 20683 8421
rect 20625 8412 20637 8415
rect 20588 8384 20637 8412
rect 20588 8372 20594 8384
rect 20625 8381 20637 8384
rect 20671 8381 20683 8415
rect 20625 8375 20683 8381
rect 20717 8415 20775 8421
rect 20717 8381 20729 8415
rect 20763 8381 20775 8415
rect 20824 8412 20852 8452
rect 21542 8440 21548 8492
rect 21600 8440 21606 8492
rect 21726 8440 21732 8492
rect 21784 8440 21790 8492
rect 21818 8440 21824 8492
rect 21876 8440 21882 8492
rect 21928 8452 22416 8480
rect 21637 8415 21695 8421
rect 21637 8412 21649 8415
rect 20824 8384 21649 8412
rect 20717 8375 20775 8381
rect 21637 8381 21649 8384
rect 21683 8412 21695 8415
rect 21928 8412 21956 8452
rect 21683 8384 21956 8412
rect 21683 8381 21695 8384
rect 21637 8375 21695 8381
rect 15120 8344 15148 8372
rect 15120 8316 15976 8344
rect 14918 8276 14924 8288
rect 14476 8248 14924 8276
rect 14918 8236 14924 8248
rect 14976 8236 14982 8288
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 15841 8279 15899 8285
rect 15841 8276 15853 8279
rect 15344 8248 15853 8276
rect 15344 8236 15350 8248
rect 15841 8245 15853 8248
rect 15887 8245 15899 8279
rect 15948 8276 15976 8316
rect 16022 8304 16028 8356
rect 16080 8344 16086 8356
rect 17402 8344 17408 8356
rect 16080 8316 17408 8344
rect 16080 8304 16086 8316
rect 17402 8304 17408 8316
rect 17460 8304 17466 8356
rect 20732 8344 20760 8375
rect 20732 8316 22048 8344
rect 22020 8288 22048 8316
rect 22094 8304 22100 8356
rect 22152 8353 22158 8356
rect 22388 8353 22416 8452
rect 22480 8421 22508 8520
rect 22465 8415 22523 8421
rect 22465 8381 22477 8415
rect 22511 8381 22523 8415
rect 22465 8375 22523 8381
rect 22152 8347 22215 8353
rect 22152 8313 22169 8347
rect 22203 8313 22215 8347
rect 22152 8307 22215 8313
rect 22373 8347 22431 8353
rect 22373 8313 22385 8347
rect 22419 8344 22431 8347
rect 22738 8344 22744 8356
rect 22419 8316 22744 8344
rect 22419 8313 22431 8316
rect 22373 8307 22431 8313
rect 22152 8304 22158 8307
rect 22738 8304 22744 8316
rect 22796 8304 22802 8356
rect 16669 8279 16727 8285
rect 16669 8276 16681 8279
rect 15948 8248 16681 8276
rect 15841 8239 15899 8245
rect 16669 8245 16681 8248
rect 16715 8276 16727 8279
rect 17195 8279 17253 8285
rect 17195 8276 17207 8279
rect 16715 8248 17207 8276
rect 16715 8245 16727 8248
rect 16669 8239 16727 8245
rect 17195 8245 17207 8248
rect 17241 8276 17253 8279
rect 17678 8276 17684 8288
rect 17241 8248 17684 8276
rect 17241 8245 17253 8248
rect 17195 8239 17253 8245
rect 17678 8236 17684 8248
rect 17736 8236 17742 8288
rect 21082 8236 21088 8288
rect 21140 8236 21146 8288
rect 22002 8236 22008 8288
rect 22060 8236 22066 8288
rect 22646 8236 22652 8288
rect 22704 8236 22710 8288
rect 552 8186 23368 8208
rect 552 8134 19022 8186
rect 19074 8134 19086 8186
rect 19138 8134 19150 8186
rect 19202 8134 19214 8186
rect 19266 8134 19278 8186
rect 19330 8134 23368 8186
rect 552 8112 23368 8134
rect 7742 8032 7748 8084
rect 7800 8032 7806 8084
rect 7837 8075 7895 8081
rect 7837 8041 7849 8075
rect 7883 8072 7895 8075
rect 8386 8072 8392 8084
rect 7883 8044 8392 8072
rect 7883 8041 7895 8044
rect 7837 8035 7895 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 10029 8075 10087 8081
rect 10029 8041 10041 8075
rect 10075 8072 10087 8075
rect 10075 8044 10824 8072
rect 10075 8041 10087 8044
rect 10029 8035 10087 8041
rect 10796 8016 10824 8044
rect 10962 8032 10968 8084
rect 11020 8032 11026 8084
rect 12526 8032 12532 8084
rect 12584 8032 12590 8084
rect 12710 8032 12716 8084
rect 12768 8032 12774 8084
rect 13170 8032 13176 8084
rect 13228 8032 13234 8084
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 13722 8072 13728 8084
rect 13320 8044 13728 8072
rect 13320 8032 13326 8044
rect 13722 8032 13728 8044
rect 13780 8072 13786 8084
rect 14182 8072 14188 8084
rect 13780 8044 14188 8072
rect 13780 8032 13786 8044
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 15749 8075 15807 8081
rect 14384 8044 15240 8072
rect 6632 8007 6690 8013
rect 6632 7973 6644 8007
rect 6678 8004 6690 8007
rect 7282 8004 7288 8016
rect 6678 7976 7288 8004
rect 6678 7973 6690 7976
rect 6632 7967 6690 7973
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 9493 8007 9551 8013
rect 8864 7976 9260 8004
rect 5902 7896 5908 7948
rect 5960 7936 5966 7948
rect 6365 7939 6423 7945
rect 6365 7936 6377 7939
rect 5960 7908 6377 7936
rect 5960 7896 5966 7908
rect 6365 7905 6377 7908
rect 6411 7936 6423 7939
rect 7098 7936 7104 7948
rect 6411 7908 7104 7936
rect 6411 7905 6423 7908
rect 6365 7899 6423 7905
rect 7098 7896 7104 7908
rect 7156 7936 7162 7948
rect 8864 7936 8892 7976
rect 7156 7908 8892 7936
rect 7156 7896 7162 7908
rect 8938 7896 8944 7948
rect 8996 7945 9002 7948
rect 9232 7945 9260 7976
rect 9493 7973 9505 8007
rect 9539 8004 9551 8007
rect 9582 8004 9588 8016
rect 9539 7976 9588 8004
rect 9539 7973 9551 7976
rect 9493 7967 9551 7973
rect 9582 7964 9588 7976
rect 9640 7964 9646 8016
rect 10229 8007 10287 8013
rect 10229 7973 10241 8007
rect 10275 8004 10287 8007
rect 10686 8004 10692 8016
rect 10275 7976 10692 8004
rect 10275 7973 10287 7976
rect 10229 7967 10287 7973
rect 10686 7964 10692 7976
rect 10744 7964 10750 8016
rect 10778 7964 10784 8016
rect 10836 7964 10842 8016
rect 12728 8004 12756 8032
rect 13050 8007 13108 8013
rect 13050 8004 13062 8007
rect 11348 7976 12480 8004
rect 12728 7976 13062 8004
rect 10778 7961 10836 7964
rect 8996 7899 9008 7945
rect 9217 7939 9275 7945
rect 9217 7905 9229 7939
rect 9263 7936 9275 7939
rect 9309 7939 9367 7945
rect 9309 7936 9321 7939
rect 9263 7908 9321 7936
rect 9263 7905 9275 7908
rect 9217 7899 9275 7905
rect 9309 7905 9321 7908
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 10152 7908 10364 7936
rect 8996 7896 9002 7899
rect 10152 7868 10180 7908
rect 9876 7840 10180 7868
rect 9876 7812 9904 7840
rect 9858 7760 9864 7812
rect 9916 7760 9922 7812
rect 10336 7800 10364 7908
rect 10502 7896 10508 7948
rect 10560 7896 10566 7948
rect 10778 7927 10790 7961
rect 10824 7927 10836 7961
rect 11348 7948 11376 7976
rect 10778 7921 10836 7927
rect 11330 7896 11336 7948
rect 11388 7896 11394 7948
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 12452 7945 12480 7976
rect 13050 7973 13062 7976
rect 13096 7973 13108 8007
rect 13188 8004 13216 8032
rect 14200 8004 14228 8032
rect 14384 8004 14412 8044
rect 13188 7976 13492 8004
rect 14200 7976 14412 8004
rect 14461 8007 14519 8013
rect 13050 7967 13108 7973
rect 12078 7939 12136 7945
rect 12078 7936 12090 7939
rect 11756 7908 12090 7936
rect 11756 7896 11762 7908
rect 12078 7905 12090 7908
rect 12124 7905 12136 7939
rect 12078 7899 12136 7905
rect 12437 7939 12495 7945
rect 12437 7905 12449 7939
rect 12483 7905 12495 7939
rect 12437 7899 12495 7905
rect 12618 7896 12624 7948
rect 12676 7936 12682 7948
rect 12713 7939 12771 7945
rect 12713 7936 12725 7939
rect 12676 7908 12725 7936
rect 12676 7896 12682 7908
rect 12713 7905 12725 7908
rect 12759 7905 12771 7939
rect 12713 7899 12771 7905
rect 12805 7939 12863 7945
rect 12805 7905 12817 7939
rect 12851 7936 12863 7939
rect 13354 7936 13360 7948
rect 12851 7908 13360 7936
rect 12851 7905 12863 7908
rect 12805 7899 12863 7905
rect 11238 7828 11244 7880
rect 11296 7828 11302 7880
rect 12345 7871 12403 7877
rect 12345 7868 12357 7871
rect 12303 7840 12357 7868
rect 12345 7837 12357 7840
rect 12391 7868 12403 7871
rect 12820 7868 12848 7899
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 13464 7936 13492 7976
rect 14461 7973 14473 8007
rect 14507 7973 14519 8007
rect 14461 7967 14519 7973
rect 14476 7936 14504 7967
rect 13464 7908 14320 7936
rect 12391 7840 12848 7868
rect 12391 7837 12403 7840
rect 12345 7831 12403 7837
rect 11256 7800 11284 7828
rect 10336 7772 11284 7800
rect 10042 7692 10048 7744
rect 10100 7692 10106 7744
rect 10318 7692 10324 7744
rect 10376 7692 10382 7744
rect 11422 7692 11428 7744
rect 11480 7732 11486 7744
rect 12360 7732 12388 7831
rect 14292 7809 14320 7908
rect 14384 7908 14504 7936
rect 14384 7868 14412 7908
rect 14734 7896 14740 7948
rect 14792 7936 14798 7948
rect 14921 7939 14979 7945
rect 14921 7936 14933 7939
rect 14792 7908 14933 7936
rect 14792 7896 14798 7908
rect 14921 7905 14933 7908
rect 14967 7905 14979 7939
rect 14921 7899 14979 7905
rect 15010 7896 15016 7948
rect 15068 7896 15074 7948
rect 15102 7896 15108 7948
rect 15160 7896 15166 7948
rect 15212 7945 15240 8044
rect 15749 8041 15761 8075
rect 15795 8072 15807 8075
rect 16022 8072 16028 8084
rect 15795 8044 16028 8072
rect 15795 8041 15807 8044
rect 15749 8035 15807 8041
rect 16022 8032 16028 8044
rect 16080 8032 16086 8084
rect 17218 8032 17224 8084
rect 17276 8072 17282 8084
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 17276 8044 17509 8072
rect 17276 8032 17282 8044
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 17497 8035 17555 8041
rect 21450 8032 21456 8084
rect 21508 8072 21514 8084
rect 21818 8072 21824 8084
rect 21508 8044 21824 8072
rect 21508 8032 21514 8044
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 22646 8072 22652 8084
rect 22572 8044 22652 8072
rect 15933 8007 15991 8013
rect 15933 7973 15945 8007
rect 15979 8004 15991 8007
rect 17865 8007 17923 8013
rect 17865 8004 17877 8007
rect 15979 7976 17877 8004
rect 15979 7973 15991 7976
rect 15933 7967 15991 7973
rect 17865 7973 17877 7976
rect 17911 7973 17923 8007
rect 17865 7967 17923 7973
rect 15197 7939 15255 7945
rect 15197 7905 15209 7939
rect 15243 7905 15255 7939
rect 15197 7899 15255 7905
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 15120 7868 15148 7896
rect 15672 7868 15700 7899
rect 16114 7896 16120 7948
rect 16172 7896 16178 7948
rect 16390 7945 16396 7948
rect 16384 7899 16396 7945
rect 16390 7896 16396 7899
rect 16448 7896 16454 7948
rect 17402 7896 17408 7948
rect 17460 7936 17466 7948
rect 17589 7939 17647 7945
rect 17589 7936 17601 7939
rect 17460 7908 17601 7936
rect 17460 7896 17466 7908
rect 17589 7905 17601 7908
rect 17635 7905 17647 7939
rect 17589 7899 17647 7905
rect 17678 7896 17684 7948
rect 17736 7896 17742 7948
rect 22572 7945 22600 8044
rect 22646 8032 22652 8044
rect 22704 8032 22710 8084
rect 22566 7939 22624 7945
rect 22566 7905 22578 7939
rect 22612 7905 22624 7939
rect 22566 7899 22624 7905
rect 22738 7896 22744 7948
rect 22796 7936 22802 7948
rect 22833 7939 22891 7945
rect 22833 7936 22845 7939
rect 22796 7908 22845 7936
rect 22796 7896 22802 7908
rect 22833 7905 22845 7908
rect 22879 7905 22891 7939
rect 22833 7899 22891 7905
rect 14384 7840 15056 7868
rect 15120 7840 15700 7868
rect 14277 7803 14335 7809
rect 14277 7769 14289 7803
rect 14323 7769 14335 7803
rect 14277 7763 14335 7769
rect 11480 7704 12388 7732
rect 11480 7692 11486 7704
rect 12710 7692 12716 7744
rect 12768 7692 12774 7744
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 14384 7732 14412 7840
rect 14826 7760 14832 7812
rect 14884 7760 14890 7812
rect 15028 7800 15056 7840
rect 17126 7828 17132 7880
rect 17184 7868 17190 7880
rect 17865 7871 17923 7877
rect 17865 7868 17877 7871
rect 17184 7840 17877 7868
rect 17184 7828 17190 7840
rect 17865 7837 17877 7840
rect 17911 7868 17923 7871
rect 19978 7868 19984 7880
rect 17911 7840 19984 7868
rect 17911 7837 17923 7840
rect 17865 7831 17923 7837
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 15102 7800 15108 7812
rect 15028 7772 15108 7800
rect 15102 7760 15108 7772
rect 15160 7760 15166 7812
rect 12860 7704 14412 7732
rect 14461 7735 14519 7741
rect 12860 7692 12866 7704
rect 14461 7701 14473 7735
rect 14507 7732 14519 7735
rect 15381 7735 15439 7741
rect 15381 7732 15393 7735
rect 14507 7704 15393 7732
rect 14507 7701 14519 7704
rect 14461 7695 14519 7701
rect 15381 7701 15393 7704
rect 15427 7701 15439 7735
rect 15381 7695 15439 7701
rect 15838 7692 15844 7744
rect 15896 7732 15902 7744
rect 15933 7735 15991 7741
rect 15933 7732 15945 7735
rect 15896 7704 15945 7732
rect 15896 7692 15902 7704
rect 15933 7701 15945 7704
rect 15979 7701 15991 7735
rect 15933 7695 15991 7701
rect 552 7642 23368 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 23368 7642
rect 552 7568 23368 7590
rect 7837 7531 7895 7537
rect 7837 7497 7849 7531
rect 7883 7528 7895 7531
rect 8202 7528 8208 7540
rect 7883 7500 8208 7528
rect 7883 7497 7895 7500
rect 7837 7491 7895 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 8757 7531 8815 7537
rect 8352 7500 8708 7528
rect 8352 7488 8358 7500
rect 5721 7463 5779 7469
rect 5721 7429 5733 7463
rect 5767 7460 5779 7463
rect 5810 7460 5816 7472
rect 5767 7432 5816 7460
rect 5767 7429 5779 7432
rect 5721 7423 5779 7429
rect 5810 7420 5816 7432
rect 5868 7420 5874 7472
rect 7653 7463 7711 7469
rect 7653 7429 7665 7463
rect 7699 7429 7711 7463
rect 7653 7423 7711 7429
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 5316 7364 7328 7392
rect 5316 7352 5322 7364
rect 5997 7259 6055 7265
rect 5997 7225 6009 7259
rect 6043 7256 6055 7259
rect 6178 7256 6184 7268
rect 6043 7228 6184 7256
rect 6043 7225 6055 7228
rect 5997 7219 6055 7225
rect 6178 7216 6184 7228
rect 6236 7216 6242 7268
rect 7300 7256 7328 7364
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 7668 7324 7696 7423
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 8481 7463 8539 7469
rect 8481 7460 8493 7463
rect 8168 7432 8493 7460
rect 8168 7420 8174 7432
rect 8220 7401 8248 7432
rect 8481 7429 8493 7432
rect 8527 7429 8539 7463
rect 8481 7423 8539 7429
rect 8680 7401 8708 7500
rect 8757 7497 8769 7531
rect 8803 7528 8815 7531
rect 8938 7528 8944 7540
rect 8803 7500 8944 7528
rect 8803 7497 8815 7500
rect 8757 7491 8815 7497
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 9769 7531 9827 7537
rect 9769 7497 9781 7531
rect 9815 7528 9827 7531
rect 10318 7528 10324 7540
rect 9815 7500 10324 7528
rect 9815 7497 9827 7500
rect 9769 7491 9827 7497
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 10502 7488 10508 7540
rect 10560 7488 10566 7540
rect 11698 7488 11704 7540
rect 11756 7488 11762 7540
rect 12526 7488 12532 7540
rect 12584 7488 12590 7540
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 12713 7531 12771 7537
rect 12713 7528 12725 7531
rect 12676 7500 12725 7528
rect 12676 7488 12682 7500
rect 12713 7497 12725 7500
rect 12759 7497 12771 7531
rect 12713 7491 12771 7497
rect 13173 7531 13231 7537
rect 13173 7497 13185 7531
rect 13219 7528 13231 7531
rect 13262 7528 13268 7540
rect 13219 7500 13268 7528
rect 13219 7497 13231 7500
rect 13173 7491 13231 7497
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 13357 7531 13415 7537
rect 13357 7497 13369 7531
rect 13403 7528 13415 7531
rect 14826 7528 14832 7540
rect 13403 7500 14832 7528
rect 13403 7497 13415 7500
rect 13357 7491 13415 7497
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 14918 7488 14924 7540
rect 14976 7488 14982 7540
rect 16945 7531 17003 7537
rect 15028 7500 16528 7528
rect 9309 7463 9367 7469
rect 9309 7429 9321 7463
rect 9355 7460 9367 7463
rect 9674 7460 9680 7472
rect 9355 7432 9680 7460
rect 9355 7429 9367 7432
rect 9309 7423 9367 7429
rect 9674 7420 9680 7432
rect 9732 7420 9738 7472
rect 9858 7420 9864 7472
rect 9916 7420 9922 7472
rect 9950 7420 9956 7472
rect 10008 7420 10014 7472
rect 10042 7420 10048 7472
rect 10100 7460 10106 7472
rect 10520 7460 10548 7488
rect 10100 7432 10548 7460
rect 12544 7460 12572 7488
rect 12544 7432 12940 7460
rect 10100 7420 10106 7432
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8665 7395 8723 7401
rect 8665 7361 8677 7395
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 9876 7392 9904 7420
rect 9447 7364 9904 7392
rect 10152 7364 10364 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 7423 7296 7696 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 8386 7284 8392 7336
rect 8444 7284 8450 7336
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7324 8999 7327
rect 9030 7324 9036 7336
rect 8987 7296 9036 7324
rect 8987 7293 8999 7296
rect 8941 7287 8999 7293
rect 7466 7256 7472 7268
rect 7300 7228 7472 7256
rect 7466 7216 7472 7228
rect 7524 7256 7530 7268
rect 7837 7259 7895 7265
rect 7837 7256 7849 7259
rect 7524 7228 7849 7256
rect 7524 7216 7530 7228
rect 7837 7225 7849 7228
rect 7883 7225 7895 7259
rect 7837 7219 7895 7225
rect 8665 7259 8723 7265
rect 8665 7225 8677 7259
rect 8711 7256 8723 7259
rect 8772 7256 8800 7287
rect 9030 7284 9036 7296
rect 9088 7284 9094 7336
rect 9125 7327 9183 7333
rect 9125 7293 9137 7327
rect 9171 7324 9183 7327
rect 10152 7324 10180 7364
rect 9171 7296 10180 7324
rect 9171 7293 9183 7296
rect 9125 7287 9183 7293
rect 10226 7284 10232 7336
rect 10284 7284 10290 7336
rect 10336 7324 10364 7364
rect 11348 7364 12572 7392
rect 11348 7336 11376 7364
rect 10686 7324 10692 7336
rect 10336 7296 10692 7324
rect 10686 7284 10692 7296
rect 10744 7284 10750 7336
rect 11330 7284 11336 7336
rect 11388 7284 11394 7336
rect 11422 7284 11428 7336
rect 11480 7284 11486 7336
rect 11532 7333 11560 7364
rect 11517 7327 11575 7333
rect 11517 7293 11529 7327
rect 11563 7293 11575 7327
rect 11517 7287 11575 7293
rect 11606 7284 11612 7336
rect 11664 7324 11670 7336
rect 11701 7327 11759 7333
rect 11701 7324 11713 7327
rect 11664 7296 11713 7324
rect 11664 7284 11670 7296
rect 11701 7293 11713 7296
rect 11747 7293 11759 7327
rect 12544 7324 12572 7364
rect 12618 7352 12624 7404
rect 12676 7352 12682 7404
rect 12912 7333 12940 7432
rect 14550 7420 14556 7472
rect 14608 7460 14614 7472
rect 15028 7460 15056 7500
rect 14608 7432 15056 7460
rect 16500 7460 16528 7500
rect 16945 7497 16957 7531
rect 16991 7528 17003 7531
rect 17402 7528 17408 7540
rect 16991 7500 17408 7528
rect 16991 7497 17003 7500
rect 16945 7491 17003 7497
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 20441 7531 20499 7537
rect 17512 7500 20392 7528
rect 17512 7460 17540 7500
rect 16500 7432 17540 7460
rect 20073 7463 20131 7469
rect 14608 7420 14614 7432
rect 20073 7429 20085 7463
rect 20119 7429 20131 7463
rect 20073 7423 20131 7429
rect 20088 7336 20116 7423
rect 20162 7420 20168 7472
rect 20220 7460 20226 7472
rect 20257 7463 20315 7469
rect 20257 7460 20269 7463
rect 20220 7432 20269 7460
rect 20220 7420 20226 7432
rect 20257 7429 20269 7432
rect 20303 7429 20315 7463
rect 20364 7460 20392 7500
rect 20441 7497 20453 7531
rect 20487 7528 20499 7531
rect 20530 7528 20536 7540
rect 20487 7500 20536 7528
rect 20487 7497 20499 7500
rect 20441 7491 20499 7497
rect 20530 7488 20536 7500
rect 20588 7488 20594 7540
rect 22097 7531 22155 7537
rect 22097 7497 22109 7531
rect 22143 7528 22155 7531
rect 22186 7528 22192 7540
rect 22143 7500 22192 7528
rect 22143 7497 22155 7500
rect 22097 7491 22155 7497
rect 22186 7488 22192 7500
rect 22244 7488 22250 7540
rect 20364 7432 22232 7460
rect 20257 7423 20315 7429
rect 21545 7395 21603 7401
rect 21545 7361 21557 7395
rect 21591 7361 21603 7395
rect 21545 7355 21603 7361
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 12544 7296 12817 7324
rect 11701 7287 11759 7293
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7324 12955 7327
rect 12943 7296 13032 7324
rect 12943 7293 12955 7296
rect 12897 7287 12955 7293
rect 8711 7228 8800 7256
rect 9309 7259 9367 7265
rect 8711 7225 8723 7228
rect 8665 7219 8723 7225
rect 9309 7225 9321 7259
rect 9355 7256 9367 7259
rect 10244 7256 10272 7284
rect 9355 7228 10272 7256
rect 9355 7225 9367 7228
rect 9309 7219 9367 7225
rect 5537 7191 5595 7197
rect 5537 7157 5549 7191
rect 5583 7188 5595 7191
rect 5626 7188 5632 7200
rect 5583 7160 5632 7188
rect 5583 7157 5595 7160
rect 5537 7151 5595 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 7558 7148 7564 7200
rect 7616 7148 7622 7200
rect 7852 7188 7880 7219
rect 11146 7216 11152 7268
rect 11204 7265 11210 7268
rect 11204 7219 11216 7265
rect 12820 7256 12848 7287
rect 13004 7268 13032 7296
rect 13354 7284 13360 7336
rect 13412 7324 13418 7336
rect 13541 7327 13599 7333
rect 13541 7324 13553 7327
rect 13412 7296 13553 7324
rect 13412 7284 13418 7296
rect 13541 7293 13553 7296
rect 13587 7324 13599 7327
rect 14366 7324 14372 7336
rect 13587 7296 14372 7324
rect 13587 7293 13599 7296
rect 13541 7287 13599 7293
rect 14366 7284 14372 7296
rect 14424 7284 14430 7336
rect 15838 7333 15844 7336
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7293 15623 7327
rect 15832 7324 15844 7333
rect 15799 7296 15844 7324
rect 15565 7287 15623 7293
rect 15832 7287 15844 7296
rect 12820 7228 12940 7256
rect 11204 7216 11210 7219
rect 9769 7191 9827 7197
rect 9769 7188 9781 7191
rect 7852 7160 9781 7188
rect 9769 7157 9781 7160
rect 9815 7188 9827 7191
rect 12802 7188 12808 7200
rect 9815 7160 12808 7188
rect 9815 7157 9827 7160
rect 9769 7151 9827 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 12912 7188 12940 7228
rect 12986 7216 12992 7268
rect 13044 7216 13050 7268
rect 13808 7259 13866 7265
rect 13808 7225 13820 7259
rect 13854 7256 13866 7259
rect 14090 7256 14096 7268
rect 13854 7228 14096 7256
rect 13854 7225 13866 7228
rect 13808 7219 13866 7225
rect 14090 7216 14096 7228
rect 14148 7216 14154 7268
rect 15580 7256 15608 7287
rect 15838 7284 15844 7287
rect 15896 7284 15902 7336
rect 16114 7284 16120 7336
rect 16172 7284 16178 7336
rect 19153 7327 19211 7333
rect 19153 7293 19165 7327
rect 19199 7324 19211 7327
rect 19518 7324 19524 7336
rect 19199 7296 19524 7324
rect 19199 7293 19211 7296
rect 19153 7287 19211 7293
rect 19518 7284 19524 7296
rect 19576 7284 19582 7336
rect 19797 7327 19855 7333
rect 19797 7293 19809 7327
rect 19843 7293 19855 7327
rect 19797 7287 19855 7293
rect 16132 7256 16160 7284
rect 19812 7256 19840 7287
rect 20070 7284 20076 7336
rect 20128 7284 20134 7336
rect 20165 7327 20223 7333
rect 20165 7293 20177 7327
rect 20211 7293 20223 7327
rect 21560 7324 21588 7355
rect 22094 7324 22100 7336
rect 21560 7296 22100 7324
rect 20165 7287 20223 7293
rect 20180 7256 20208 7287
rect 22094 7284 22100 7296
rect 22152 7284 22158 7336
rect 22204 7333 22232 7432
rect 22189 7327 22247 7333
rect 22189 7293 22201 7327
rect 22235 7324 22247 7327
rect 22278 7324 22284 7336
rect 22235 7296 22284 7324
rect 22235 7293 22247 7296
rect 22189 7287 22247 7293
rect 22278 7284 22284 7296
rect 22336 7284 22342 7336
rect 22465 7327 22523 7333
rect 22465 7293 22477 7327
rect 22511 7324 22523 7327
rect 22830 7324 22836 7336
rect 22511 7296 22836 7324
rect 22511 7293 22523 7296
rect 22465 7287 22523 7293
rect 22830 7284 22836 7296
rect 22888 7284 22894 7336
rect 20625 7259 20683 7265
rect 20625 7256 20637 7259
rect 15580 7228 16160 7256
rect 19444 7228 20116 7256
rect 20180 7228 20637 7256
rect 19444 7200 19472 7228
rect 13189 7191 13247 7197
rect 13189 7188 13201 7191
rect 12912 7160 13201 7188
rect 13189 7157 13201 7160
rect 13235 7188 13247 7191
rect 14734 7188 14740 7200
rect 13235 7160 14740 7188
rect 13235 7157 13247 7160
rect 13189 7151 13247 7157
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 18414 7148 18420 7200
rect 18472 7188 18478 7200
rect 19061 7191 19119 7197
rect 19061 7188 19073 7191
rect 18472 7160 19073 7188
rect 18472 7148 18478 7160
rect 19061 7157 19073 7160
rect 19107 7157 19119 7191
rect 19061 7151 19119 7157
rect 19426 7148 19432 7200
rect 19484 7148 19490 7200
rect 19794 7148 19800 7200
rect 19852 7188 19858 7200
rect 19889 7191 19947 7197
rect 19889 7188 19901 7191
rect 19852 7160 19901 7188
rect 19852 7148 19858 7160
rect 19889 7157 19901 7160
rect 19935 7157 19947 7191
rect 19889 7151 19947 7157
rect 19978 7148 19984 7200
rect 20036 7148 20042 7200
rect 20088 7188 20116 7228
rect 20625 7225 20637 7228
rect 20671 7256 20683 7259
rect 20714 7256 20720 7268
rect 20671 7228 20720 7256
rect 20671 7225 20683 7228
rect 20625 7219 20683 7225
rect 20714 7216 20720 7228
rect 20772 7216 20778 7268
rect 21729 7259 21787 7265
rect 21729 7225 21741 7259
rect 21775 7256 21787 7259
rect 22554 7256 22560 7268
rect 21775 7228 22560 7256
rect 21775 7225 21787 7228
rect 21729 7219 21787 7225
rect 22554 7216 22560 7228
rect 22612 7216 22618 7268
rect 20415 7191 20473 7197
rect 20415 7188 20427 7191
rect 20088 7160 20427 7188
rect 20415 7157 20427 7160
rect 20461 7157 20473 7191
rect 20415 7151 20473 7157
rect 21634 7148 21640 7200
rect 21692 7148 21698 7200
rect 552 7098 23368 7120
rect 552 7046 19022 7098
rect 19074 7046 19086 7098
rect 19138 7046 19150 7098
rect 19202 7046 19214 7098
rect 19266 7046 19278 7098
rect 19330 7046 23368 7098
rect 552 7024 23368 7046
rect 4724 6956 5396 6984
rect 4724 6780 4752 6956
rect 5261 6919 5319 6925
rect 5261 6885 5273 6919
rect 5307 6885 5319 6919
rect 5261 6879 5319 6885
rect 4801 6851 4859 6857
rect 4801 6817 4813 6851
rect 4847 6848 4859 6851
rect 4847 6820 5120 6848
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 4264 6752 4752 6780
rect 4264 6656 4292 6752
rect 5092 6721 5120 6820
rect 5276 6780 5304 6879
rect 5368 6848 5396 6956
rect 9950 6944 9956 6996
rect 10008 6944 10014 6996
rect 10686 6944 10692 6996
rect 10744 6984 10750 6996
rect 10781 6987 10839 6993
rect 10781 6984 10793 6987
rect 10744 6956 10793 6984
rect 10744 6944 10750 6956
rect 10781 6953 10793 6956
rect 10827 6953 10839 6987
rect 10781 6947 10839 6953
rect 11146 6944 11152 6996
rect 11204 6944 11210 6996
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 12768 6956 12848 6984
rect 12768 6944 12774 6956
rect 6178 6876 6184 6928
rect 6236 6916 6242 6928
rect 6549 6919 6607 6925
rect 6549 6916 6561 6919
rect 6236 6888 6561 6916
rect 6236 6876 6242 6888
rect 6549 6885 6561 6888
rect 6595 6885 6607 6919
rect 6549 6879 6607 6885
rect 7558 6876 7564 6928
rect 7616 6916 7622 6928
rect 9674 6925 9680 6928
rect 7714 6919 7772 6925
rect 7714 6916 7726 6919
rect 7616 6888 7726 6916
rect 7616 6876 7622 6888
rect 7714 6885 7726 6888
rect 7760 6885 7772 6919
rect 7714 6879 7772 6885
rect 9668 6879 9680 6925
rect 9674 6876 9680 6879
rect 9732 6876 9738 6928
rect 6089 6851 6147 6857
rect 6089 6848 6101 6851
rect 5368 6820 6101 6848
rect 6089 6817 6101 6820
rect 6135 6848 6147 6851
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 6135 6820 6469 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 6457 6817 6469 6820
rect 6503 6817 6515 6851
rect 6733 6851 6791 6857
rect 6733 6848 6745 6851
rect 6457 6811 6515 6817
rect 6656 6820 6745 6848
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5276 6752 5825 6780
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 5902 6740 5908 6792
rect 5960 6780 5966 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5960 6752 6009 6780
rect 5960 6740 5966 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 5077 6715 5135 6721
rect 5077 6681 5089 6715
rect 5123 6681 5135 6715
rect 5077 6675 5135 6681
rect 5350 6672 5356 6724
rect 5408 6712 5414 6724
rect 5629 6715 5687 6721
rect 5629 6712 5641 6715
rect 5408 6684 5641 6712
rect 5408 6672 5414 6684
rect 5629 6681 5641 6684
rect 5675 6681 5687 6715
rect 6012 6712 6040 6743
rect 6178 6740 6184 6792
rect 6236 6740 6242 6792
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 6472 6780 6500 6811
rect 6546 6780 6552 6792
rect 6472 6752 6552 6780
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 6656 6712 6684 6820
rect 6733 6817 6745 6820
rect 6779 6817 6791 6851
rect 6733 6811 6791 6817
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 7469 6851 7527 6857
rect 7469 6848 7481 6851
rect 7156 6820 7481 6848
rect 7156 6808 7162 6820
rect 7469 6817 7481 6820
rect 7515 6817 7527 6851
rect 9968 6848 9996 6944
rect 12820 6925 12848 6956
rect 12986 6944 12992 6996
rect 13044 6984 13050 6996
rect 13909 6987 13967 6993
rect 13909 6984 13921 6987
rect 13044 6956 13921 6984
rect 13044 6944 13050 6956
rect 13909 6953 13921 6956
rect 13955 6953 13967 6987
rect 13909 6947 13967 6953
rect 12796 6919 12854 6925
rect 12796 6885 12808 6919
rect 12842 6885 12854 6919
rect 13924 6916 13952 6947
rect 14090 6944 14096 6996
rect 14148 6944 14154 6996
rect 16301 6987 16359 6993
rect 16301 6953 16313 6987
rect 16347 6984 16359 6987
rect 16390 6984 16396 6996
rect 16347 6956 16396 6984
rect 16347 6953 16359 6956
rect 16301 6947 16359 6953
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 18138 6944 18144 6996
rect 18196 6984 18202 6996
rect 18575 6987 18633 6993
rect 18575 6984 18587 6987
rect 18196 6956 18587 6984
rect 18196 6944 18202 6956
rect 18575 6953 18587 6956
rect 18621 6953 18633 6987
rect 19702 6984 19708 6996
rect 18575 6947 18633 6953
rect 18800 6956 19708 6984
rect 15010 6916 15016 6928
rect 13924 6888 15016 6916
rect 12796 6879 12854 6885
rect 15010 6876 15016 6888
rect 15068 6876 15074 6928
rect 15286 6876 15292 6928
rect 15344 6916 15350 6928
rect 18800 6925 18828 6956
rect 19702 6944 19708 6956
rect 19760 6984 19766 6996
rect 20070 6984 20076 6996
rect 19760 6956 20076 6984
rect 19760 6944 19766 6956
rect 20070 6944 20076 6956
rect 20128 6944 20134 6996
rect 20438 6944 20444 6996
rect 20496 6944 20502 6996
rect 20714 6944 20720 6996
rect 20772 6984 20778 6996
rect 21358 6984 21364 6996
rect 20772 6956 21364 6984
rect 20772 6944 20778 6956
rect 21358 6944 21364 6956
rect 21416 6944 21422 6996
rect 21634 6944 21640 6996
rect 21692 6984 21698 6996
rect 21729 6987 21787 6993
rect 21729 6984 21741 6987
rect 21692 6956 21741 6984
rect 21692 6944 21698 6956
rect 21729 6953 21741 6956
rect 21775 6953 21787 6987
rect 21729 6947 21787 6953
rect 22281 6987 22339 6993
rect 22281 6953 22293 6987
rect 22327 6953 22339 6987
rect 22281 6947 22339 6953
rect 18785 6919 18843 6925
rect 18785 6916 18797 6919
rect 15344 6888 18797 6916
rect 15344 6876 15350 6888
rect 18785 6885 18797 6888
rect 18831 6885 18843 6919
rect 18785 6879 18843 6885
rect 19978 6876 19984 6928
rect 20036 6876 20042 6928
rect 20254 6876 20260 6928
rect 20312 6876 20318 6928
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 9968 6820 10977 6848
rect 7469 6811 7527 6817
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 10965 6811 11023 6817
rect 13998 6808 14004 6860
rect 14056 6808 14062 6860
rect 14185 6851 14243 6857
rect 14185 6817 14197 6851
rect 14231 6848 14243 6851
rect 14642 6848 14648 6860
rect 14231 6820 14648 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 15654 6808 15660 6860
rect 15712 6848 15718 6860
rect 16117 6851 16175 6857
rect 16117 6848 16129 6851
rect 15712 6820 16129 6848
rect 15712 6808 15718 6820
rect 16117 6817 16129 6820
rect 16163 6817 16175 6851
rect 16117 6811 16175 6817
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6848 18199 6851
rect 18187 6820 18460 6848
rect 18187 6817 18199 6820
rect 18141 6811 18199 6817
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6749 9459 6783
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 9401 6743 9459 6749
rect 12406 6752 12541 6780
rect 7006 6712 7012 6724
rect 6012 6684 6684 6712
rect 6748 6684 7012 6712
rect 5629 6675 5687 6681
rect 4246 6604 4252 6656
rect 4304 6604 4310 6656
rect 4985 6647 5043 6653
rect 4985 6613 4997 6647
rect 5031 6644 5043 6647
rect 5166 6644 5172 6656
rect 5031 6616 5172 6644
rect 5031 6613 5043 6616
rect 4985 6607 5043 6613
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 5258 6604 5264 6656
rect 5316 6604 5322 6656
rect 5644 6644 5672 6675
rect 6748 6644 6776 6684
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 5644 6616 6776 6644
rect 6914 6604 6920 6656
rect 6972 6604 6978 6656
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 8849 6647 8907 6653
rect 8849 6644 8861 6647
rect 8628 6616 8861 6644
rect 8628 6604 8634 6616
rect 8849 6613 8861 6616
rect 8895 6613 8907 6647
rect 9416 6644 9444 6743
rect 11422 6644 11428 6656
rect 9416 6616 11428 6644
rect 8849 6607 8907 6613
rect 11422 6604 11428 6616
rect 11480 6644 11486 6656
rect 12406 6644 12434 6752
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 18432 6721 18460 6820
rect 18874 6808 18880 6860
rect 18932 6848 18938 6860
rect 19061 6851 19119 6857
rect 19061 6848 19073 6851
rect 18932 6820 19073 6848
rect 18932 6808 18938 6820
rect 19061 6817 19073 6820
rect 19107 6817 19119 6851
rect 19061 6811 19119 6817
rect 19076 6780 19104 6811
rect 19150 6808 19156 6860
rect 19208 6848 19214 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 19208 6820 19257 6848
rect 19208 6808 19214 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 19613 6851 19671 6857
rect 19613 6817 19625 6851
rect 19659 6817 19671 6851
rect 19613 6811 19671 6817
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 19076 6752 19441 6780
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 18417 6715 18475 6721
rect 18417 6681 18429 6715
rect 18463 6681 18475 6715
rect 18417 6675 18475 6681
rect 18782 6672 18788 6724
rect 18840 6712 18846 6724
rect 19150 6712 19156 6724
rect 18840 6684 19156 6712
rect 18840 6672 18846 6684
rect 19150 6672 19156 6684
rect 19208 6672 19214 6724
rect 19444 6712 19472 6743
rect 19518 6740 19524 6792
rect 19576 6780 19582 6792
rect 19628 6780 19656 6811
rect 19886 6808 19892 6860
rect 19944 6808 19950 6860
rect 19996 6848 20024 6876
rect 20346 6848 20352 6860
rect 19996 6820 20352 6848
rect 20346 6808 20352 6820
rect 20404 6848 20410 6860
rect 20732 6857 20760 6944
rect 21082 6876 21088 6928
rect 21140 6916 21146 6928
rect 21140 6888 22048 6916
rect 21140 6876 21146 6888
rect 22020 6860 22048 6888
rect 22186 6876 22192 6928
rect 22244 6916 22250 6928
rect 22296 6916 22324 6947
rect 22554 6944 22560 6996
rect 22612 6944 22618 6996
rect 22738 6944 22744 6996
rect 22796 6944 22802 6996
rect 22756 6916 22784 6944
rect 22244 6888 22784 6916
rect 22244 6876 22250 6888
rect 20533 6851 20591 6857
rect 20533 6848 20545 6851
rect 20404 6820 20545 6848
rect 20404 6808 20410 6820
rect 20533 6817 20545 6820
rect 20579 6817 20591 6851
rect 20533 6811 20591 6817
rect 20717 6851 20775 6857
rect 20717 6817 20729 6851
rect 20763 6817 20775 6851
rect 20717 6811 20775 6817
rect 20809 6851 20867 6857
rect 20809 6817 20821 6851
rect 20855 6848 20867 6851
rect 20898 6848 20904 6860
rect 20855 6820 20904 6848
rect 20855 6817 20867 6820
rect 20809 6811 20867 6817
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 21361 6851 21419 6857
rect 21361 6848 21373 6851
rect 21008 6820 21373 6848
rect 19576 6772 20576 6780
rect 20622 6772 20628 6792
rect 19576 6752 20628 6772
rect 19576 6740 19582 6752
rect 20548 6744 20628 6752
rect 20622 6740 20628 6744
rect 20680 6740 20686 6792
rect 19702 6712 19708 6724
rect 19444 6684 19708 6712
rect 19702 6672 19708 6684
rect 19760 6672 19766 6724
rect 20806 6672 20812 6724
rect 20864 6672 20870 6724
rect 21008 6721 21036 6820
rect 21361 6817 21373 6820
rect 21407 6817 21419 6851
rect 21361 6811 21419 6817
rect 22002 6808 22008 6860
rect 22060 6808 22066 6860
rect 22097 6851 22155 6857
rect 22097 6817 22109 6851
rect 22143 6817 22155 6851
rect 22097 6811 22155 6817
rect 21450 6740 21456 6792
rect 21508 6740 21514 6792
rect 21821 6783 21879 6789
rect 21821 6780 21833 6783
rect 21560 6752 21833 6780
rect 20993 6715 21051 6721
rect 20993 6681 21005 6715
rect 21039 6681 21051 6715
rect 21560 6712 21588 6752
rect 21821 6749 21833 6752
rect 21867 6780 21879 6783
rect 21910 6780 21916 6792
rect 21867 6752 21916 6780
rect 21867 6749 21879 6752
rect 21821 6743 21879 6749
rect 21910 6740 21916 6752
rect 21968 6740 21974 6792
rect 22112 6712 22140 6811
rect 22462 6808 22468 6860
rect 22520 6808 22526 6860
rect 22557 6851 22615 6857
rect 22557 6817 22569 6851
rect 22603 6848 22615 6851
rect 22603 6820 22692 6848
rect 22603 6817 22615 6820
rect 22557 6811 22615 6817
rect 20993 6675 21051 6681
rect 21468 6684 21588 6712
rect 21836 6684 22140 6712
rect 11480 6616 12434 6644
rect 11480 6604 11486 6616
rect 18322 6604 18328 6656
rect 18380 6604 18386 6656
rect 18601 6647 18659 6653
rect 18601 6613 18613 6647
rect 18647 6644 18659 6647
rect 18877 6647 18935 6653
rect 18877 6644 18889 6647
rect 18647 6616 18889 6644
rect 18647 6613 18659 6616
rect 18601 6607 18659 6613
rect 18877 6613 18889 6616
rect 18923 6613 18935 6647
rect 18877 6607 18935 6613
rect 19794 6604 19800 6656
rect 19852 6604 19858 6656
rect 20070 6604 20076 6656
rect 20128 6644 20134 6656
rect 20257 6647 20315 6653
rect 20257 6644 20269 6647
rect 20128 6616 20269 6644
rect 20128 6604 20134 6616
rect 20257 6613 20269 6616
rect 20303 6613 20315 6647
rect 20257 6607 20315 6613
rect 20622 6604 20628 6656
rect 20680 6604 20686 6656
rect 20824 6644 20852 6672
rect 21468 6644 21496 6684
rect 20824 6616 21496 6644
rect 21542 6604 21548 6656
rect 21600 6644 21606 6656
rect 21836 6644 21864 6684
rect 21600 6616 21864 6644
rect 21600 6604 21606 6616
rect 21910 6604 21916 6656
rect 21968 6604 21974 6656
rect 22094 6604 22100 6656
rect 22152 6644 22158 6656
rect 22664 6644 22692 6820
rect 22738 6808 22744 6860
rect 22796 6808 22802 6860
rect 22152 6616 22692 6644
rect 22152 6604 22158 6616
rect 552 6554 23368 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 23368 6554
rect 552 6480 23368 6502
rect 6178 6440 6184 6452
rect 4816 6412 6184 6440
rect 4816 6304 4844 6412
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 6328 6412 6377 6440
rect 6328 6400 6334 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 4816 6276 4936 6304
rect 4338 6196 4344 6248
rect 4396 6196 4402 6248
rect 4908 6245 4936 6276
rect 4801 6239 4859 6245
rect 4801 6236 4813 6239
rect 4540 6208 4813 6236
rect 4540 6168 4568 6208
rect 4801 6205 4813 6208
rect 4847 6205 4859 6239
rect 4801 6199 4859 6205
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 4985 6239 5043 6245
rect 4985 6205 4997 6239
rect 5031 6236 5043 6239
rect 5074 6236 5080 6248
rect 5031 6208 5080 6236
rect 5031 6205 5043 6208
rect 4985 6199 5043 6205
rect 5074 6196 5080 6208
rect 5132 6196 5138 6248
rect 5258 6245 5264 6248
rect 5241 6239 5264 6245
rect 5241 6205 5253 6239
rect 5241 6199 5264 6205
rect 5258 6196 5264 6199
rect 5316 6196 5322 6248
rect 6380 6236 6408 6403
rect 7006 6400 7012 6452
rect 7064 6400 7070 6452
rect 18322 6400 18328 6452
rect 18380 6400 18386 6452
rect 18874 6400 18880 6452
rect 18932 6440 18938 6452
rect 20073 6443 20131 6449
rect 20073 6440 20085 6443
rect 18932 6412 20085 6440
rect 18932 6400 18938 6412
rect 20073 6409 20085 6412
rect 20119 6409 20131 6443
rect 20073 6403 20131 6409
rect 20254 6400 20260 6452
rect 20312 6440 20318 6452
rect 20901 6443 20959 6449
rect 20901 6440 20913 6443
rect 20312 6412 20913 6440
rect 20312 6400 20318 6412
rect 20901 6409 20913 6412
rect 20947 6409 20959 6443
rect 22738 6440 22744 6452
rect 20901 6403 20959 6409
rect 21192 6412 21680 6440
rect 17604 6344 18184 6372
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 6880 6276 7328 6304
rect 6880 6264 6886 6276
rect 7300 6245 7328 6276
rect 7650 6264 7656 6316
rect 7708 6264 7714 6316
rect 17604 6245 17632 6344
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6304 17739 6307
rect 17727 6276 18092 6304
rect 17727 6273 17739 6276
rect 17681 6267 17739 6273
rect 6733 6239 6791 6245
rect 6733 6236 6745 6239
rect 6380 6208 6745 6236
rect 6733 6205 6745 6208
rect 6779 6205 6791 6239
rect 6733 6199 6791 6205
rect 7193 6239 7251 6245
rect 7193 6205 7205 6239
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 17589 6239 17647 6245
rect 17589 6205 17601 6239
rect 17635 6205 17647 6239
rect 17589 6199 17647 6205
rect 17773 6239 17831 6245
rect 17773 6205 17785 6239
rect 17819 6205 17831 6239
rect 17773 6199 17831 6205
rect 4264 6140 4568 6168
rect 4617 6171 4675 6177
rect 4264 6112 4292 6140
rect 4617 6137 4629 6171
rect 4663 6168 4675 6171
rect 5902 6168 5908 6180
rect 4663 6140 5908 6168
rect 4663 6137 4675 6140
rect 4617 6131 4675 6137
rect 5902 6128 5908 6140
rect 5960 6128 5966 6180
rect 6270 6128 6276 6180
rect 6328 6168 6334 6180
rect 6457 6171 6515 6177
rect 6457 6168 6469 6171
rect 6328 6140 6469 6168
rect 6328 6128 6334 6140
rect 6457 6137 6469 6140
rect 6503 6137 6515 6171
rect 6825 6171 6883 6177
rect 6825 6168 6837 6171
rect 6457 6131 6515 6137
rect 6564 6140 6837 6168
rect 4246 6060 4252 6112
rect 4304 6060 4310 6112
rect 4522 6060 4528 6112
rect 4580 6060 4586 6112
rect 4890 6060 4896 6112
rect 4948 6060 4954 6112
rect 5920 6100 5948 6128
rect 6362 6100 6368 6112
rect 5920 6072 6368 6100
rect 6362 6060 6368 6072
rect 6420 6100 6426 6112
rect 6564 6100 6592 6140
rect 6825 6137 6837 6140
rect 6871 6137 6883 6171
rect 6825 6131 6883 6137
rect 6420 6072 6592 6100
rect 6420 6060 6426 6072
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 7208 6100 7236 6199
rect 17788 6168 17816 6199
rect 17862 6196 17868 6248
rect 17920 6196 17926 6248
rect 18064 6245 18092 6276
rect 18156 6248 18184 6344
rect 18340 6304 18368 6400
rect 19794 6332 19800 6384
rect 19852 6372 19858 6384
rect 20530 6372 20536 6384
rect 19852 6344 20536 6372
rect 19852 6332 19858 6344
rect 20530 6332 20536 6344
rect 20588 6372 20594 6384
rect 21192 6372 21220 6412
rect 20588 6344 21220 6372
rect 20588 6332 20594 6344
rect 18340 6276 18828 6304
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 18138 6196 18144 6248
rect 18196 6196 18202 6248
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6236 18291 6239
rect 18414 6236 18420 6248
rect 18279 6208 18420 6236
rect 18279 6205 18291 6208
rect 18233 6199 18291 6205
rect 18248 6168 18276 6199
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 18690 6196 18696 6248
rect 18748 6196 18754 6248
rect 18800 6236 18828 6276
rect 20180 6276 20668 6304
rect 20180 6248 20208 6276
rect 18949 6239 19007 6245
rect 18949 6236 18961 6239
rect 18800 6208 18961 6236
rect 18949 6205 18961 6208
rect 18995 6205 19007 6239
rect 18949 6199 19007 6205
rect 19886 6196 19892 6248
rect 19944 6196 19950 6248
rect 20162 6196 20168 6248
rect 20220 6196 20226 6248
rect 20346 6196 20352 6248
rect 20404 6236 20410 6248
rect 20640 6245 20668 6276
rect 21082 6264 21088 6316
rect 21140 6264 21146 6316
rect 21192 6313 21220 6344
rect 21450 6332 21456 6384
rect 21508 6372 21514 6384
rect 21545 6375 21603 6381
rect 21545 6372 21557 6375
rect 21508 6344 21557 6372
rect 21508 6332 21514 6344
rect 21545 6341 21557 6344
rect 21591 6341 21603 6375
rect 21652 6372 21680 6412
rect 22066 6412 22744 6440
rect 22066 6372 22094 6412
rect 22738 6400 22744 6412
rect 22796 6400 22802 6452
rect 21652 6344 22094 6372
rect 21545 6335 21603 6341
rect 22646 6332 22652 6384
rect 22704 6332 22710 6384
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6273 21235 6307
rect 21177 6267 21235 6273
rect 22002 6264 22008 6316
rect 22060 6304 22066 6316
rect 22060 6276 22416 6304
rect 22060 6264 22066 6276
rect 20441 6239 20499 6245
rect 20441 6236 20453 6239
rect 20404 6208 20453 6236
rect 20404 6196 20410 6208
rect 20441 6205 20453 6208
rect 20487 6205 20499 6239
rect 20441 6199 20499 6205
rect 20533 6239 20591 6245
rect 20533 6205 20545 6239
rect 20579 6205 20591 6239
rect 20533 6199 20591 6205
rect 20625 6239 20683 6245
rect 20625 6205 20637 6239
rect 20671 6205 20683 6239
rect 20625 6199 20683 6205
rect 17788 6140 18276 6168
rect 19904 6168 19932 6196
rect 20548 6168 20576 6199
rect 20806 6196 20812 6248
rect 20864 6196 20870 6248
rect 21269 6239 21327 6245
rect 21269 6205 21281 6239
rect 21315 6205 21327 6239
rect 21269 6199 21327 6205
rect 19904 6140 20576 6168
rect 21284 6168 21312 6199
rect 21358 6196 21364 6248
rect 21416 6196 21422 6248
rect 21818 6196 21824 6248
rect 21876 6236 21882 6248
rect 22388 6245 22416 6276
rect 21913 6239 21971 6245
rect 21913 6236 21925 6239
rect 21876 6208 21925 6236
rect 21876 6196 21882 6208
rect 21913 6205 21925 6208
rect 21959 6205 21971 6239
rect 22373 6239 22431 6245
rect 21913 6199 21971 6205
rect 22020 6208 22232 6236
rect 21542 6168 21548 6180
rect 21284 6140 21548 6168
rect 21542 6128 21548 6140
rect 21600 6168 21606 6180
rect 21729 6171 21787 6177
rect 21729 6168 21741 6171
rect 21600 6140 21741 6168
rect 21600 6128 21606 6140
rect 21729 6137 21741 6140
rect 21775 6168 21787 6171
rect 22020 6168 22048 6208
rect 21775 6140 22048 6168
rect 21775 6137 21787 6140
rect 21729 6131 21787 6137
rect 22094 6128 22100 6180
rect 22152 6128 22158 6180
rect 22204 6168 22232 6208
rect 22373 6205 22385 6239
rect 22419 6205 22431 6239
rect 22373 6199 22431 6205
rect 22554 6196 22560 6248
rect 22612 6196 22618 6248
rect 22830 6196 22836 6248
rect 22888 6196 22894 6248
rect 22572 6168 22600 6196
rect 22204 6140 22600 6168
rect 6696 6072 7236 6100
rect 6696 6060 6702 6072
rect 7374 6060 7380 6112
rect 7432 6060 7438 6112
rect 18506 6060 18512 6112
rect 18564 6060 18570 6112
rect 20162 6060 20168 6112
rect 20220 6060 20226 6112
rect 21358 6060 21364 6112
rect 21416 6100 21422 6112
rect 21821 6103 21879 6109
rect 21821 6100 21833 6103
rect 21416 6072 21833 6100
rect 21416 6060 21422 6072
rect 21821 6069 21833 6072
rect 21867 6069 21879 6103
rect 21821 6063 21879 6069
rect 22002 6060 22008 6112
rect 22060 6100 22066 6112
rect 22189 6103 22247 6109
rect 22189 6100 22201 6103
rect 22060 6072 22201 6100
rect 22060 6060 22066 6072
rect 22189 6069 22201 6072
rect 22235 6069 22247 6103
rect 22189 6063 22247 6069
rect 552 6010 23368 6032
rect 552 5958 19022 6010
rect 19074 5958 19086 6010
rect 19138 5958 19150 6010
rect 19202 5958 19214 6010
rect 19266 5958 19278 6010
rect 19330 5958 23368 6010
rect 552 5936 23368 5958
rect 4246 5856 4252 5908
rect 4304 5856 4310 5908
rect 4338 5856 4344 5908
rect 4396 5856 4402 5908
rect 4890 5856 4896 5908
rect 4948 5856 4954 5908
rect 5074 5856 5080 5908
rect 5132 5896 5138 5908
rect 5810 5896 5816 5908
rect 5132 5868 5816 5896
rect 5132 5856 5138 5868
rect 5810 5856 5816 5868
rect 5868 5856 5874 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7443 5899 7501 5905
rect 7443 5896 7455 5899
rect 6972 5868 7455 5896
rect 6972 5856 6978 5868
rect 7443 5865 7455 5868
rect 7489 5865 7501 5899
rect 7443 5859 7501 5865
rect 18506 5856 18512 5908
rect 18564 5856 18570 5908
rect 19429 5899 19487 5905
rect 19429 5865 19441 5899
rect 19475 5896 19487 5899
rect 19518 5896 19524 5908
rect 19475 5868 19524 5896
rect 19475 5865 19487 5868
rect 19429 5859 19487 5865
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 20162 5856 20168 5908
rect 20220 5856 20226 5908
rect 20346 5856 20352 5908
rect 20404 5896 20410 5908
rect 21085 5899 21143 5905
rect 21085 5896 21097 5899
rect 20404 5868 21097 5896
rect 20404 5856 20410 5868
rect 21085 5865 21097 5868
rect 21131 5896 21143 5899
rect 21818 5896 21824 5908
rect 21131 5868 21824 5896
rect 21131 5865 21143 5868
rect 21085 5859 21143 5865
rect 21818 5856 21824 5868
rect 21876 5856 21882 5908
rect 22554 5856 22560 5908
rect 22612 5896 22618 5908
rect 22833 5899 22891 5905
rect 22833 5896 22845 5899
rect 22612 5868 22845 5896
rect 22612 5856 22618 5868
rect 22833 5865 22845 5868
rect 22879 5865 22891 5899
rect 22833 5859 22891 5865
rect 4356 5556 4384 5856
rect 4908 5828 4936 5856
rect 7653 5831 7711 5837
rect 7653 5828 7665 5831
rect 4908 5800 7665 5828
rect 7653 5797 7665 5800
rect 7699 5797 7711 5831
rect 7653 5791 7711 5797
rect 18316 5831 18374 5837
rect 18316 5797 18328 5831
rect 18362 5828 18374 5831
rect 18524 5828 18552 5856
rect 18362 5800 18552 5828
rect 19972 5831 20030 5837
rect 18362 5797 18374 5800
rect 18316 5791 18374 5797
rect 19972 5797 19984 5831
rect 20018 5828 20030 5831
rect 20180 5828 20208 5856
rect 22186 5828 22192 5840
rect 20018 5800 20208 5828
rect 21468 5800 22192 5828
rect 20018 5797 20030 5800
rect 19972 5791 20030 5797
rect 5373 5763 5431 5769
rect 5373 5729 5385 5763
rect 5419 5760 5431 5763
rect 5534 5760 5540 5772
rect 5419 5732 5540 5760
rect 5419 5729 5431 5732
rect 5373 5723 5431 5729
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5729 5687 5763
rect 5629 5723 5687 5729
rect 5644 5692 5672 5723
rect 5718 5720 5724 5772
rect 5776 5760 5782 5772
rect 6069 5763 6127 5769
rect 6069 5760 6081 5763
rect 5776 5732 6081 5760
rect 5776 5720 5782 5732
rect 6069 5729 6081 5732
rect 6115 5729 6127 5763
rect 6069 5723 6127 5729
rect 18049 5763 18107 5769
rect 18049 5729 18061 5763
rect 18095 5760 18107 5763
rect 18690 5760 18696 5772
rect 18095 5732 18696 5760
rect 18095 5729 18107 5732
rect 18049 5723 18107 5729
rect 18690 5720 18696 5732
rect 18748 5760 18754 5772
rect 19705 5763 19763 5769
rect 19705 5760 19717 5763
rect 18748 5732 19717 5760
rect 18748 5720 18754 5732
rect 19705 5729 19717 5732
rect 19751 5760 19763 5763
rect 19794 5760 19800 5772
rect 19751 5732 19800 5760
rect 19751 5729 19763 5732
rect 19705 5723 19763 5729
rect 19794 5720 19800 5732
rect 19852 5760 19858 5772
rect 21468 5769 21496 5800
rect 22186 5788 22192 5800
rect 22244 5788 22250 5840
rect 21726 5769 21732 5772
rect 21453 5763 21511 5769
rect 21453 5760 21465 5763
rect 19852 5732 21465 5760
rect 19852 5720 19858 5732
rect 21453 5729 21465 5732
rect 21499 5729 21511 5763
rect 21453 5723 21511 5729
rect 21720 5723 21732 5769
rect 21726 5720 21732 5723
rect 21784 5720 21790 5772
rect 5810 5692 5816 5704
rect 5644 5664 5816 5692
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 7285 5627 7343 5633
rect 7285 5624 7297 5627
rect 6748 5596 7297 5624
rect 6748 5556 6776 5596
rect 7285 5593 7297 5596
rect 7331 5593 7343 5627
rect 7285 5587 7343 5593
rect 4356 5528 6776 5556
rect 6822 5516 6828 5568
rect 6880 5556 6886 5568
rect 7193 5559 7251 5565
rect 7193 5556 7205 5559
rect 6880 5528 7205 5556
rect 6880 5516 6886 5528
rect 7193 5525 7205 5528
rect 7239 5525 7251 5559
rect 7193 5519 7251 5525
rect 7466 5516 7472 5568
rect 7524 5516 7530 5568
rect 552 5466 23368 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 23368 5466
rect 552 5392 23368 5414
rect 4985 5355 5043 5361
rect 4985 5321 4997 5355
rect 5031 5352 5043 5355
rect 5718 5352 5724 5364
rect 5031 5324 5724 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 6362 5312 6368 5364
rect 6420 5352 6426 5364
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 6420 5324 6469 5352
rect 6420 5312 6426 5324
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 18877 5355 18935 5361
rect 18877 5352 18889 5355
rect 18196 5324 18889 5352
rect 18196 5312 18202 5324
rect 18877 5321 18889 5324
rect 18923 5321 18935 5355
rect 18877 5315 18935 5321
rect 21358 5312 21364 5364
rect 21416 5312 21422 5364
rect 21637 5355 21695 5361
rect 21637 5321 21649 5355
rect 21683 5352 21695 5355
rect 21726 5352 21732 5364
rect 21683 5324 21732 5352
rect 21683 5321 21695 5324
rect 21637 5315 21695 5321
rect 21726 5312 21732 5324
rect 21784 5312 21790 5364
rect 4816 5188 5212 5216
rect 4522 5108 4528 5160
rect 4580 5108 4586 5160
rect 4816 5157 4844 5188
rect 4801 5151 4859 5157
rect 4801 5117 4813 5151
rect 4847 5117 4859 5151
rect 4801 5111 4859 5117
rect 5074 5108 5080 5160
rect 5132 5108 5138 5160
rect 5184 5148 5212 5188
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6822 5216 6828 5228
rect 6328 5188 6828 5216
rect 6328 5176 6334 5188
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 19794 5176 19800 5228
rect 19852 5216 19858 5228
rect 19981 5219 20039 5225
rect 19981 5216 19993 5219
rect 19852 5188 19993 5216
rect 19852 5176 19858 5188
rect 19981 5185 19993 5188
rect 20027 5185 20039 5219
rect 22002 5216 22008 5228
rect 19981 5179 20039 5185
rect 21468 5188 22008 5216
rect 5626 5148 5632 5160
rect 5184 5120 5632 5148
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 18782 5108 18788 5160
rect 18840 5108 18846 5160
rect 18874 5108 18880 5160
rect 18932 5148 18938 5160
rect 21468 5157 21496 5188
rect 22002 5176 22008 5188
rect 22060 5176 22066 5228
rect 18969 5151 19027 5157
rect 18969 5148 18981 5151
rect 18932 5120 18981 5148
rect 18932 5108 18938 5120
rect 18969 5117 18981 5120
rect 19015 5117 19027 5151
rect 21453 5151 21511 5157
rect 21453 5148 21465 5151
rect 18969 5111 19027 5117
rect 20180 5120 21465 5148
rect 4540 5080 4568 5108
rect 5322 5083 5380 5089
rect 5322 5080 5334 5083
rect 4540 5052 5334 5080
rect 5322 5049 5334 5052
rect 5368 5049 5380 5083
rect 18800 5080 18828 5108
rect 20180 5080 20208 5120
rect 21453 5117 21465 5120
rect 21499 5117 21511 5151
rect 21453 5111 21511 5117
rect 21637 5151 21695 5157
rect 21637 5117 21649 5151
rect 21683 5148 21695 5151
rect 21910 5148 21916 5160
rect 21683 5120 21916 5148
rect 21683 5117 21695 5120
rect 21637 5111 21695 5117
rect 21910 5108 21916 5120
rect 21968 5108 21974 5160
rect 20254 5089 20260 5092
rect 18800 5052 20208 5080
rect 5322 5043 5380 5049
rect 20248 5043 20260 5089
rect 20254 5040 20260 5043
rect 20312 5040 20318 5092
rect 552 4922 23368 4944
rect 552 4870 19022 4922
rect 19074 4870 19086 4922
rect 19138 4870 19150 4922
rect 19202 4870 19214 4922
rect 19266 4870 19278 4922
rect 19330 4870 23368 4922
rect 552 4848 23368 4870
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5813 4811 5871 4817
rect 5813 4808 5825 4811
rect 5592 4780 5825 4808
rect 5592 4768 5598 4780
rect 5813 4777 5825 4780
rect 5859 4777 5871 4811
rect 5813 4771 5871 4777
rect 20254 4768 20260 4820
rect 20312 4768 20318 4820
rect 20438 4768 20444 4820
rect 20496 4768 20502 4820
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 7374 4672 7380 4684
rect 6043 4644 7380 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 20456 4681 20484 4768
rect 20441 4675 20499 4681
rect 20441 4641 20453 4675
rect 20487 4641 20499 4675
rect 20441 4635 20499 4641
rect 6270 4564 6276 4616
rect 6328 4564 6334 4616
rect 6638 4564 6644 4616
rect 6696 4564 6702 4616
rect 6181 4539 6239 4545
rect 6181 4505 6193 4539
rect 6227 4536 6239 4539
rect 6656 4536 6684 4564
rect 6227 4508 6684 4536
rect 6227 4505 6239 4508
rect 6181 4499 6239 4505
rect 552 4378 23368 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 23368 4378
rect 552 4304 23368 4326
rect 22278 4088 22284 4140
rect 22336 4128 22342 4140
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 22336 4100 22753 4128
rect 22336 4088 22342 4100
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 22741 4091 22799 4097
rect 23014 4020 23020 4072
rect 23072 4020 23078 4072
rect 552 3834 23368 3856
rect 552 3782 19022 3834
rect 19074 3782 19086 3834
rect 19138 3782 19150 3834
rect 19202 3782 19214 3834
rect 19266 3782 19278 3834
rect 19330 3782 23368 3834
rect 552 3760 23368 3782
rect 552 3290 23368 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 23368 3290
rect 552 3216 23368 3238
rect 552 2746 23368 2768
rect 552 2694 19022 2746
rect 19074 2694 19086 2746
rect 19138 2694 19150 2746
rect 19202 2694 19214 2746
rect 19266 2694 19278 2746
rect 19330 2694 23368 2746
rect 552 2672 23368 2694
rect 552 2202 23368 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 23368 2202
rect 552 2128 23368 2150
rect 552 1658 23368 1680
rect 552 1606 19022 1658
rect 19074 1606 19086 1658
rect 19138 1606 19150 1658
rect 19202 1606 19214 1658
rect 19266 1606 19278 1658
rect 19330 1606 23368 1658
rect 552 1584 23368 1606
rect 552 1114 23368 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 23368 1114
rect 552 1040 23368 1062
rect 552 570 23368 592
rect 552 518 19022 570
rect 19074 518 19086 570
rect 19138 518 19150 570
rect 19202 518 19214 570
rect 19266 518 19278 570
rect 19330 518 23368 570
rect 552 496 23368 518
<< via1 >>
rect 15936 23468 15988 23520
rect 18420 23468 18472 23520
rect 19022 23366 19074 23418
rect 19086 23366 19138 23418
rect 19150 23366 19202 23418
rect 19214 23366 19266 23418
rect 19278 23366 19330 23418
rect 1676 23264 1728 23316
rect 11520 23264 11572 23316
rect 4620 23196 4672 23248
rect 7564 23196 7616 23248
rect 5816 23171 5868 23180
rect 5816 23137 5825 23171
rect 5825 23137 5859 23171
rect 5859 23137 5868 23171
rect 5816 23128 5868 23137
rect 7196 23128 7248 23180
rect 7656 23128 7708 23180
rect 5908 23060 5960 23112
rect 9680 23103 9732 23112
rect 9680 23069 9689 23103
rect 9689 23069 9723 23103
rect 9723 23069 9732 23103
rect 9680 23060 9732 23069
rect 4344 22924 4396 22976
rect 4896 22967 4948 22976
rect 4896 22933 4905 22967
rect 4905 22933 4939 22967
rect 4939 22933 4948 22967
rect 4896 22924 4948 22933
rect 6644 22992 6696 23044
rect 10140 22992 10192 23044
rect 7104 22967 7156 22976
rect 7104 22933 7113 22967
rect 7113 22933 7147 22967
rect 7147 22933 7156 22967
rect 7104 22924 7156 22933
rect 7472 22924 7524 22976
rect 9496 22924 9548 22976
rect 10324 23103 10376 23112
rect 10324 23069 10333 23103
rect 10333 23069 10367 23103
rect 10367 23069 10376 23103
rect 10324 23060 10376 23069
rect 10692 23196 10744 23248
rect 14372 23196 14424 23248
rect 10508 23171 10560 23180
rect 10508 23137 10517 23171
rect 10517 23137 10551 23171
rect 10551 23137 10560 23171
rect 10508 23128 10560 23137
rect 13452 23128 13504 23180
rect 15200 23196 15252 23248
rect 15936 23171 15988 23180
rect 15936 23137 15945 23171
rect 15945 23137 15979 23171
rect 15979 23137 15988 23171
rect 15936 23128 15988 23137
rect 20904 23264 20956 23316
rect 17040 23196 17092 23248
rect 11796 23103 11848 23112
rect 11796 23069 11805 23103
rect 11805 23069 11839 23103
rect 11839 23069 11848 23103
rect 11796 23060 11848 23069
rect 14556 23060 14608 23112
rect 14924 22992 14976 23044
rect 11244 22924 11296 22976
rect 14648 22924 14700 22976
rect 16304 23103 16356 23112
rect 16304 23069 16313 23103
rect 16313 23069 16347 23103
rect 16347 23069 16356 23103
rect 16304 23060 16356 23069
rect 17040 22992 17092 23044
rect 16120 22924 16172 22976
rect 17500 23128 17552 23180
rect 18696 23171 18748 23180
rect 18696 23137 18705 23171
rect 18705 23137 18739 23171
rect 18739 23137 18748 23171
rect 18696 23128 18748 23137
rect 19340 23128 19392 23180
rect 19432 23171 19484 23180
rect 19432 23137 19441 23171
rect 19441 23137 19475 23171
rect 19475 23137 19484 23171
rect 19432 23128 19484 23137
rect 20536 23196 20588 23248
rect 20720 23171 20772 23180
rect 18420 23060 18472 23112
rect 19892 23060 19944 23112
rect 20720 23137 20729 23171
rect 20729 23137 20763 23171
rect 20763 23137 20772 23171
rect 20720 23128 20772 23137
rect 22284 23128 22336 23180
rect 17776 22924 17828 22976
rect 19064 22924 19116 22976
rect 19616 22924 19668 22976
rect 20996 23060 21048 23112
rect 21548 22924 21600 22976
rect 3662 22822 3714 22874
rect 3726 22822 3778 22874
rect 3790 22822 3842 22874
rect 3854 22822 3906 22874
rect 3918 22822 3970 22874
rect 5816 22720 5868 22772
rect 5264 22652 5316 22704
rect 4620 22516 4672 22568
rect 4896 22516 4948 22568
rect 5908 22559 5960 22568
rect 5908 22525 5917 22559
rect 5917 22525 5951 22559
rect 5951 22525 5960 22559
rect 5908 22516 5960 22525
rect 6184 22516 6236 22568
rect 6644 22559 6696 22568
rect 6644 22525 6655 22559
rect 6655 22525 6689 22559
rect 6689 22525 6696 22559
rect 6644 22516 6696 22525
rect 7380 22720 7432 22772
rect 7656 22720 7708 22772
rect 7196 22652 7248 22704
rect 4896 22423 4948 22432
rect 4896 22389 4905 22423
rect 4905 22389 4939 22423
rect 4939 22389 4948 22423
rect 4896 22380 4948 22389
rect 6644 22423 6696 22432
rect 6644 22389 6653 22423
rect 6653 22389 6687 22423
rect 6687 22389 6696 22423
rect 6644 22380 6696 22389
rect 7196 22448 7248 22500
rect 7472 22448 7524 22500
rect 8484 22720 8536 22772
rect 9680 22763 9732 22772
rect 9680 22729 9689 22763
rect 9689 22729 9723 22763
rect 9723 22729 9732 22763
rect 9680 22720 9732 22729
rect 10140 22720 10192 22772
rect 10324 22652 10376 22704
rect 16304 22720 16356 22772
rect 18696 22720 18748 22772
rect 8116 22627 8168 22636
rect 8116 22593 8125 22627
rect 8125 22593 8159 22627
rect 8159 22593 8168 22627
rect 8116 22584 8168 22593
rect 7932 22559 7984 22568
rect 7932 22525 7941 22559
rect 7941 22525 7975 22559
rect 7975 22525 7984 22559
rect 7932 22516 7984 22525
rect 9036 22559 9088 22568
rect 9036 22525 9045 22559
rect 9045 22525 9079 22559
rect 9079 22525 9088 22559
rect 9036 22516 9088 22525
rect 9496 22559 9548 22568
rect 9496 22525 9505 22559
rect 9505 22525 9539 22559
rect 9539 22525 9548 22559
rect 9496 22516 9548 22525
rect 10140 22516 10192 22568
rect 11428 22584 11480 22636
rect 11336 22559 11388 22568
rect 11336 22525 11345 22559
rect 11345 22525 11379 22559
rect 11379 22525 11388 22559
rect 11336 22516 11388 22525
rect 11980 22584 12032 22636
rect 8024 22448 8076 22500
rect 14372 22516 14424 22568
rect 13912 22448 13964 22500
rect 9496 22380 9548 22432
rect 12440 22380 12492 22432
rect 12532 22423 12584 22432
rect 12532 22389 12541 22423
rect 12541 22389 12575 22423
rect 12575 22389 12584 22423
rect 12532 22380 12584 22389
rect 12900 22423 12952 22432
rect 12900 22389 12909 22423
rect 12909 22389 12943 22423
rect 12943 22389 12952 22423
rect 12900 22380 12952 22389
rect 14556 22380 14608 22432
rect 14924 22516 14976 22568
rect 15384 22516 15436 22568
rect 15568 22559 15620 22568
rect 15568 22525 15577 22559
rect 15577 22525 15611 22559
rect 15611 22525 15620 22559
rect 15568 22516 15620 22525
rect 15016 22448 15068 22500
rect 17316 22516 17368 22568
rect 17408 22559 17460 22568
rect 17408 22525 17417 22559
rect 17417 22525 17451 22559
rect 17451 22525 17460 22559
rect 17408 22516 17460 22525
rect 17776 22559 17828 22568
rect 17776 22525 17785 22559
rect 17785 22525 17819 22559
rect 17819 22525 17828 22559
rect 17776 22516 17828 22525
rect 18420 22584 18472 22636
rect 19340 22584 19392 22636
rect 16580 22448 16632 22500
rect 19064 22559 19116 22568
rect 19064 22525 19073 22559
rect 19073 22525 19107 22559
rect 19107 22525 19116 22559
rect 19064 22516 19116 22525
rect 19524 22559 19576 22568
rect 19524 22525 19533 22559
rect 19533 22525 19567 22559
rect 19567 22525 19576 22559
rect 19524 22516 19576 22525
rect 19892 22559 19944 22568
rect 19892 22525 19901 22559
rect 19901 22525 19935 22559
rect 19935 22525 19944 22559
rect 19892 22516 19944 22525
rect 20996 22627 21048 22636
rect 20996 22593 21005 22627
rect 21005 22593 21039 22627
rect 21039 22593 21048 22627
rect 20996 22584 21048 22593
rect 21456 22627 21508 22636
rect 21456 22593 21465 22627
rect 21465 22593 21499 22627
rect 21499 22593 21508 22627
rect 21456 22584 21508 22593
rect 21916 22627 21968 22636
rect 21916 22593 21925 22627
rect 21925 22593 21959 22627
rect 21959 22593 21968 22627
rect 21916 22584 21968 22593
rect 15568 22380 15620 22432
rect 17500 22380 17552 22432
rect 17776 22380 17828 22432
rect 18604 22448 18656 22500
rect 21548 22559 21600 22568
rect 21548 22525 21557 22559
rect 21557 22525 21591 22559
rect 21591 22525 21600 22559
rect 21548 22516 21600 22525
rect 22008 22559 22060 22568
rect 22008 22525 22017 22559
rect 22017 22525 22051 22559
rect 22051 22525 22060 22559
rect 22008 22516 22060 22525
rect 22192 22559 22244 22568
rect 22192 22525 22201 22559
rect 22201 22525 22235 22559
rect 22235 22525 22244 22559
rect 22192 22516 22244 22525
rect 20720 22448 20772 22500
rect 19892 22380 19944 22432
rect 21088 22380 21140 22432
rect 22100 22423 22152 22432
rect 22100 22389 22109 22423
rect 22109 22389 22143 22423
rect 22143 22389 22152 22423
rect 22100 22380 22152 22389
rect 19022 22278 19074 22330
rect 19086 22278 19138 22330
rect 19150 22278 19202 22330
rect 19214 22278 19266 22330
rect 19278 22278 19330 22330
rect 4896 22176 4948 22228
rect 4344 22108 4396 22160
rect 8024 22176 8076 22228
rect 9036 22176 9088 22228
rect 9956 22176 10008 22228
rect 10508 22176 10560 22228
rect 6736 22151 6788 22160
rect 6736 22117 6745 22151
rect 6745 22117 6779 22151
rect 6779 22117 6788 22151
rect 6736 22108 6788 22117
rect 7472 22108 7524 22160
rect 7840 22108 7892 22160
rect 6460 21972 6512 22024
rect 5172 21836 5224 21888
rect 6368 21836 6420 21888
rect 6460 21879 6512 21888
rect 6460 21845 6469 21879
rect 6469 21845 6503 21879
rect 6503 21845 6512 21879
rect 6460 21836 6512 21845
rect 6828 21904 6880 21956
rect 7748 22083 7800 22092
rect 7748 22049 7757 22083
rect 7757 22049 7791 22083
rect 7791 22049 7800 22083
rect 7748 22040 7800 22049
rect 9220 22040 9272 22092
rect 9772 22040 9824 22092
rect 8484 21972 8536 22024
rect 9956 22083 10008 22092
rect 9956 22049 9965 22083
rect 9965 22049 9999 22083
rect 9999 22049 10008 22083
rect 9956 22040 10008 22049
rect 7288 21904 7340 21956
rect 7840 21904 7892 21956
rect 10140 22015 10192 22024
rect 10140 21981 10149 22015
rect 10149 21981 10183 22015
rect 10183 21981 10192 22015
rect 10140 21972 10192 21981
rect 11336 22108 11388 22160
rect 11980 22176 12032 22228
rect 11520 22040 11572 22092
rect 11704 22083 11756 22092
rect 11704 22049 11713 22083
rect 11713 22049 11747 22083
rect 11747 22049 11756 22083
rect 11704 22040 11756 22049
rect 13084 22151 13136 22160
rect 13084 22117 13093 22151
rect 13093 22117 13127 22151
rect 13127 22117 13136 22151
rect 13084 22108 13136 22117
rect 17868 22176 17920 22228
rect 18604 22176 18656 22228
rect 20996 22176 21048 22228
rect 15016 22108 15068 22160
rect 17592 22151 17644 22160
rect 17592 22117 17601 22151
rect 17601 22117 17635 22151
rect 17635 22117 17644 22151
rect 17592 22108 17644 22117
rect 10508 21947 10560 21956
rect 10508 21913 10517 21947
rect 10517 21913 10551 21947
rect 10551 21913 10560 21947
rect 10508 21904 10560 21913
rect 11428 21947 11480 21956
rect 11428 21913 11437 21947
rect 11437 21913 11471 21947
rect 11471 21913 11480 21947
rect 11428 21904 11480 21913
rect 7196 21836 7248 21888
rect 8116 21836 8168 21888
rect 8208 21879 8260 21888
rect 8208 21845 8217 21879
rect 8217 21845 8251 21879
rect 8251 21845 8260 21879
rect 8208 21836 8260 21845
rect 14464 22083 14516 22092
rect 14464 22049 14473 22083
rect 14473 22049 14507 22083
rect 14507 22049 14516 22083
rect 14464 22040 14516 22049
rect 14648 22040 14700 22092
rect 16120 22083 16172 22092
rect 16120 22049 16129 22083
rect 16129 22049 16163 22083
rect 16163 22049 16172 22083
rect 16120 22040 16172 22049
rect 17040 22040 17092 22092
rect 17500 22083 17552 22092
rect 17500 22049 17509 22083
rect 17509 22049 17543 22083
rect 17543 22049 17552 22083
rect 17500 22040 17552 22049
rect 19616 22108 19668 22160
rect 19984 22151 20036 22160
rect 19984 22117 19993 22151
rect 19993 22117 20027 22151
rect 20027 22117 20036 22151
rect 19984 22108 20036 22117
rect 14280 21972 14332 22024
rect 17868 21972 17920 22024
rect 18696 22040 18748 22092
rect 18788 22040 18840 22092
rect 19432 22083 19484 22092
rect 19432 22049 19441 22083
rect 19441 22049 19475 22083
rect 19475 22049 19484 22083
rect 19432 22040 19484 22049
rect 19524 22040 19576 22092
rect 19708 22040 19760 22092
rect 20536 22108 20588 22160
rect 20168 22083 20220 22092
rect 20168 22049 20177 22083
rect 20177 22049 20211 22083
rect 20211 22049 20220 22083
rect 20168 22040 20220 22049
rect 20260 22040 20312 22092
rect 20720 22040 20772 22092
rect 21456 22083 21508 22092
rect 21456 22049 21465 22083
rect 21465 22049 21499 22083
rect 21499 22049 21508 22083
rect 21456 22040 21508 22049
rect 22008 22176 22060 22228
rect 22192 22176 22244 22228
rect 19340 21972 19392 22024
rect 20628 21972 20680 22024
rect 20812 21972 20864 22024
rect 21916 21972 21968 22024
rect 20260 21904 20312 21956
rect 12716 21836 12768 21888
rect 14740 21836 14792 21888
rect 16948 21836 17000 21888
rect 17132 21836 17184 21888
rect 17408 21879 17460 21888
rect 17408 21845 17417 21879
rect 17417 21845 17451 21879
rect 17451 21845 17460 21879
rect 17408 21836 17460 21845
rect 18144 21879 18196 21888
rect 18144 21845 18153 21879
rect 18153 21845 18187 21879
rect 18187 21845 18196 21879
rect 18144 21836 18196 21845
rect 19432 21836 19484 21888
rect 20720 21879 20772 21888
rect 20720 21845 20729 21879
rect 20729 21845 20763 21879
rect 20763 21845 20772 21879
rect 20720 21836 20772 21845
rect 21088 21836 21140 21888
rect 3662 21734 3714 21786
rect 3726 21734 3778 21786
rect 3790 21734 3842 21786
rect 3854 21734 3906 21786
rect 3918 21734 3970 21786
rect 6828 21675 6880 21684
rect 6828 21641 6837 21675
rect 6837 21641 6871 21675
rect 6871 21641 6880 21675
rect 6828 21632 6880 21641
rect 7288 21632 7340 21684
rect 7748 21632 7800 21684
rect 9680 21632 9732 21684
rect 7656 21564 7708 21616
rect 7932 21564 7984 21616
rect 7196 21428 7248 21480
rect 7380 21428 7432 21480
rect 7748 21496 7800 21548
rect 10048 21564 10100 21616
rect 6828 21360 6880 21412
rect 9496 21428 9548 21480
rect 10232 21564 10284 21616
rect 13912 21632 13964 21684
rect 17132 21675 17184 21684
rect 17132 21641 17141 21675
rect 17141 21641 17175 21675
rect 17175 21641 17184 21675
rect 17132 21632 17184 21641
rect 8024 21360 8076 21412
rect 8760 21360 8812 21412
rect 9772 21360 9824 21412
rect 11152 21471 11204 21480
rect 11152 21437 11161 21471
rect 11161 21437 11195 21471
rect 11195 21437 11204 21471
rect 11152 21428 11204 21437
rect 12440 21539 12492 21548
rect 12440 21505 12449 21539
rect 12449 21505 12483 21539
rect 12483 21505 12492 21539
rect 12440 21496 12492 21505
rect 12532 21496 12584 21548
rect 14280 21564 14332 21616
rect 10416 21403 10468 21412
rect 10416 21369 10425 21403
rect 10425 21369 10459 21403
rect 10459 21369 10468 21403
rect 10416 21360 10468 21369
rect 10968 21360 11020 21412
rect 13820 21471 13872 21480
rect 13820 21437 13829 21471
rect 13829 21437 13863 21471
rect 13863 21437 13872 21471
rect 13820 21428 13872 21437
rect 13912 21428 13964 21480
rect 16948 21564 17000 21616
rect 19432 21632 19484 21684
rect 14740 21539 14792 21548
rect 14740 21505 14749 21539
rect 14749 21505 14783 21539
rect 14783 21505 14792 21539
rect 14740 21496 14792 21505
rect 17776 21564 17828 21616
rect 6184 21292 6236 21344
rect 7472 21292 7524 21344
rect 10876 21335 10928 21344
rect 10876 21301 10885 21335
rect 10885 21301 10919 21335
rect 10919 21301 10928 21335
rect 10876 21292 10928 21301
rect 12716 21292 12768 21344
rect 13268 21292 13320 21344
rect 14004 21403 14056 21412
rect 14004 21369 14013 21403
rect 14013 21369 14047 21403
rect 14047 21369 14056 21403
rect 14004 21360 14056 21369
rect 14648 21360 14700 21412
rect 15568 21428 15620 21480
rect 16580 21428 16632 21480
rect 16488 21360 16540 21412
rect 17592 21471 17644 21480
rect 17592 21437 17601 21471
rect 17601 21437 17635 21471
rect 17635 21437 17644 21471
rect 17592 21428 17644 21437
rect 18144 21564 18196 21616
rect 20168 21632 20220 21684
rect 20996 21632 21048 21684
rect 21272 21632 21324 21684
rect 19984 21564 20036 21616
rect 18696 21539 18748 21548
rect 18696 21505 18705 21539
rect 18705 21505 18739 21539
rect 18739 21505 18748 21539
rect 18696 21496 18748 21505
rect 18788 21428 18840 21480
rect 14280 21335 14332 21344
rect 14280 21301 14289 21335
rect 14289 21301 14323 21335
rect 14323 21301 14332 21335
rect 14280 21292 14332 21301
rect 14924 21292 14976 21344
rect 15752 21292 15804 21344
rect 16672 21292 16724 21344
rect 17868 21360 17920 21412
rect 19340 21403 19392 21412
rect 19340 21369 19349 21403
rect 19349 21369 19383 21403
rect 19383 21369 19392 21403
rect 19340 21360 19392 21369
rect 19524 21403 19576 21412
rect 19524 21369 19565 21403
rect 19565 21369 19576 21403
rect 19800 21471 19852 21480
rect 19800 21437 19809 21471
rect 19809 21437 19843 21471
rect 19843 21437 19852 21471
rect 19800 21428 19852 21437
rect 20536 21496 20588 21548
rect 20904 21496 20956 21548
rect 19524 21360 19576 21369
rect 20260 21360 20312 21412
rect 20536 21360 20588 21412
rect 20812 21360 20864 21412
rect 20996 21428 21048 21480
rect 22100 21539 22152 21548
rect 22100 21505 22109 21539
rect 22109 21505 22143 21539
rect 22143 21505 22152 21539
rect 22100 21496 22152 21505
rect 18236 21335 18288 21344
rect 18236 21301 18245 21335
rect 18245 21301 18279 21335
rect 18279 21301 18288 21335
rect 18236 21292 18288 21301
rect 21180 21292 21232 21344
rect 22008 21335 22060 21344
rect 22008 21301 22017 21335
rect 22017 21301 22051 21335
rect 22051 21301 22060 21335
rect 22008 21292 22060 21301
rect 22560 21335 22612 21344
rect 22560 21301 22569 21335
rect 22569 21301 22603 21335
rect 22603 21301 22612 21335
rect 22560 21292 22612 21301
rect 19022 21190 19074 21242
rect 19086 21190 19138 21242
rect 19150 21190 19202 21242
rect 19214 21190 19266 21242
rect 19278 21190 19330 21242
rect 6368 21088 6420 21140
rect 7288 21088 7340 21140
rect 7380 21088 7432 21140
rect 5356 21020 5408 21072
rect 4620 20952 4672 21004
rect 5632 20995 5684 21004
rect 5632 20961 5641 20995
rect 5641 20961 5675 20995
rect 5675 20961 5684 20995
rect 5632 20952 5684 20961
rect 4436 20927 4488 20936
rect 4436 20893 4445 20927
rect 4445 20893 4479 20927
rect 4479 20893 4488 20927
rect 4436 20884 4488 20893
rect 5356 20884 5408 20936
rect 6000 20995 6052 21004
rect 6000 20961 6009 20995
rect 6009 20961 6043 20995
rect 6043 20961 6052 20995
rect 6000 20952 6052 20961
rect 5264 20816 5316 20868
rect 6276 20952 6328 21004
rect 6368 20952 6420 21004
rect 7472 20952 7524 21004
rect 6828 20884 6880 20936
rect 7932 20995 7984 21004
rect 7932 20961 7941 20995
rect 7941 20961 7975 20995
rect 7975 20961 7984 20995
rect 7932 20952 7984 20961
rect 7656 20927 7708 20936
rect 7656 20893 7665 20927
rect 7665 20893 7699 20927
rect 7699 20893 7708 20927
rect 8208 21088 8260 21140
rect 10416 21088 10468 21140
rect 10876 21088 10928 21140
rect 11152 21088 11204 21140
rect 8116 20952 8168 21004
rect 10232 20952 10284 21004
rect 10968 20995 11020 21004
rect 10968 20961 10977 20995
rect 10977 20961 11011 20995
rect 11011 20961 11020 20995
rect 10968 20952 11020 20961
rect 13912 21088 13964 21140
rect 16304 21088 16356 21140
rect 11704 21020 11756 21072
rect 12808 20952 12860 21004
rect 7656 20884 7708 20893
rect 11888 20884 11940 20936
rect 13360 21020 13412 21072
rect 14648 21020 14700 21072
rect 19800 21088 19852 21140
rect 19984 21088 20036 21140
rect 14004 20952 14056 21004
rect 15200 20952 15252 21004
rect 15384 20952 15436 21004
rect 16488 20952 16540 21004
rect 16580 20952 16632 21004
rect 19708 21020 19760 21072
rect 8024 20816 8076 20868
rect 8116 20859 8168 20868
rect 8116 20825 8125 20859
rect 8125 20825 8159 20859
rect 8159 20825 8168 20859
rect 8116 20816 8168 20825
rect 12716 20859 12768 20868
rect 12716 20825 12725 20859
rect 12725 20825 12759 20859
rect 12759 20825 12768 20859
rect 12716 20816 12768 20825
rect 13452 20859 13504 20868
rect 13452 20825 13461 20859
rect 13461 20825 13495 20859
rect 13495 20825 13504 20859
rect 13452 20816 13504 20825
rect 15752 20884 15804 20936
rect 16672 20884 16724 20936
rect 17592 20952 17644 21004
rect 17960 20952 18012 21004
rect 21180 21020 21232 21072
rect 21088 20952 21140 21004
rect 21272 20995 21324 21004
rect 21272 20961 21281 20995
rect 21281 20961 21315 20995
rect 21315 20961 21324 20995
rect 21272 20952 21324 20961
rect 14464 20816 14516 20868
rect 17408 20816 17460 20868
rect 20720 20816 20772 20868
rect 21272 20816 21324 20868
rect 5172 20748 5224 20800
rect 5632 20791 5684 20800
rect 5632 20757 5641 20791
rect 5641 20757 5675 20791
rect 5675 20757 5684 20791
rect 5632 20748 5684 20757
rect 7748 20791 7800 20800
rect 7748 20757 7757 20791
rect 7757 20757 7791 20791
rect 7791 20757 7800 20791
rect 7748 20748 7800 20757
rect 11612 20748 11664 20800
rect 14556 20748 14608 20800
rect 17500 20791 17552 20800
rect 17500 20757 17509 20791
rect 17509 20757 17543 20791
rect 17543 20757 17552 20791
rect 17500 20748 17552 20757
rect 20812 20748 20864 20800
rect 21916 20791 21968 20800
rect 21916 20757 21925 20791
rect 21925 20757 21959 20791
rect 21959 20757 21968 20791
rect 21916 20748 21968 20757
rect 3662 20646 3714 20698
rect 3726 20646 3778 20698
rect 3790 20646 3842 20698
rect 3854 20646 3906 20698
rect 3918 20646 3970 20698
rect 5632 20544 5684 20596
rect 6000 20587 6052 20596
rect 6000 20553 6009 20587
rect 6009 20553 6043 20587
rect 6043 20553 6052 20587
rect 6000 20544 6052 20553
rect 7748 20544 7800 20596
rect 7932 20544 7984 20596
rect 12808 20544 12860 20596
rect 15200 20544 15252 20596
rect 18052 20544 18104 20596
rect 5816 20476 5868 20528
rect 7288 20519 7340 20528
rect 7288 20485 7297 20519
rect 7297 20485 7331 20519
rect 7331 20485 7340 20519
rect 7288 20476 7340 20485
rect 8208 20408 8260 20460
rect 4344 20383 4396 20392
rect 4344 20349 4353 20383
rect 4353 20349 4387 20383
rect 4387 20349 4396 20383
rect 4344 20340 4396 20349
rect 4436 20383 4488 20392
rect 4436 20349 4445 20383
rect 4445 20349 4479 20383
rect 4479 20349 4488 20383
rect 4436 20340 4488 20349
rect 4620 20383 4672 20392
rect 4620 20349 4629 20383
rect 4629 20349 4663 20383
rect 4663 20349 4672 20383
rect 4620 20340 4672 20349
rect 4252 20272 4304 20324
rect 5172 20383 5224 20392
rect 5172 20349 5181 20383
rect 5181 20349 5215 20383
rect 5215 20349 5224 20383
rect 5172 20340 5224 20349
rect 5264 20383 5316 20392
rect 5264 20349 5273 20383
rect 5273 20349 5307 20383
rect 5307 20349 5316 20383
rect 5264 20340 5316 20349
rect 5356 20383 5408 20392
rect 5356 20349 5365 20383
rect 5365 20349 5399 20383
rect 5399 20349 5408 20383
rect 5356 20340 5408 20349
rect 6368 20340 6420 20392
rect 7656 20340 7708 20392
rect 7932 20340 7984 20392
rect 12164 20340 12216 20392
rect 13452 20408 13504 20460
rect 12992 20340 13044 20392
rect 7104 20272 7156 20324
rect 5724 20247 5776 20256
rect 5724 20213 5733 20247
rect 5733 20213 5767 20247
rect 5767 20213 5776 20247
rect 5724 20204 5776 20213
rect 9404 20272 9456 20324
rect 8392 20204 8444 20256
rect 13360 20340 13412 20392
rect 13544 20315 13596 20324
rect 13544 20281 13553 20315
rect 13553 20281 13587 20315
rect 13587 20281 13596 20315
rect 13544 20272 13596 20281
rect 14004 20340 14056 20392
rect 14464 20383 14516 20392
rect 14464 20349 14473 20383
rect 14473 20349 14507 20383
rect 14507 20349 14516 20383
rect 14464 20340 14516 20349
rect 14556 20340 14608 20392
rect 14648 20383 14700 20392
rect 14648 20349 14657 20383
rect 14657 20349 14691 20383
rect 14691 20349 14700 20383
rect 14648 20340 14700 20349
rect 15384 20340 15436 20392
rect 17408 20340 17460 20392
rect 17500 20340 17552 20392
rect 17592 20383 17644 20392
rect 17592 20349 17601 20383
rect 17601 20349 17635 20383
rect 17635 20349 17644 20383
rect 17592 20340 17644 20349
rect 17960 20383 18012 20392
rect 17960 20349 17969 20383
rect 17969 20349 18003 20383
rect 18003 20349 18012 20383
rect 17960 20340 18012 20349
rect 18236 20340 18288 20392
rect 20812 20340 20864 20392
rect 21916 20544 21968 20596
rect 22008 20476 22060 20528
rect 21916 20408 21968 20460
rect 13728 20204 13780 20256
rect 15200 20315 15252 20324
rect 15200 20281 15209 20315
rect 15209 20281 15243 20315
rect 15243 20281 15252 20315
rect 15200 20272 15252 20281
rect 22560 20383 22612 20392
rect 22560 20349 22569 20383
rect 22569 20349 22603 20383
rect 22603 20349 22612 20383
rect 22560 20340 22612 20349
rect 16304 20204 16356 20256
rect 17224 20247 17276 20256
rect 17224 20213 17233 20247
rect 17233 20213 17267 20247
rect 17267 20213 17276 20247
rect 17224 20204 17276 20213
rect 18604 20204 18656 20256
rect 20812 20204 20864 20256
rect 21180 20247 21232 20256
rect 21180 20213 21189 20247
rect 21189 20213 21223 20247
rect 21223 20213 21232 20247
rect 21180 20204 21232 20213
rect 21456 20204 21508 20256
rect 22284 20247 22336 20256
rect 22284 20213 22293 20247
rect 22293 20213 22327 20247
rect 22327 20213 22336 20247
rect 22284 20204 22336 20213
rect 19022 20102 19074 20154
rect 19086 20102 19138 20154
rect 19150 20102 19202 20154
rect 19214 20102 19266 20154
rect 19278 20102 19330 20154
rect 5264 20000 5316 20052
rect 5356 20000 5408 20052
rect 10048 20000 10100 20052
rect 10232 19932 10284 19984
rect 11336 19932 11388 19984
rect 13084 20043 13136 20052
rect 13084 20009 13093 20043
rect 13093 20009 13127 20043
rect 13127 20009 13136 20043
rect 13084 20000 13136 20009
rect 13544 20000 13596 20052
rect 17224 20000 17276 20052
rect 17500 20000 17552 20052
rect 5724 19864 5776 19916
rect 6828 19907 6880 19916
rect 6828 19873 6837 19907
rect 6837 19873 6871 19907
rect 6871 19873 6880 19907
rect 6828 19864 6880 19873
rect 7748 19864 7800 19916
rect 8760 19907 8812 19916
rect 8760 19873 8769 19907
rect 8769 19873 8803 19907
rect 8803 19873 8812 19907
rect 8760 19864 8812 19873
rect 10048 19907 10100 19916
rect 10048 19873 10057 19907
rect 10057 19873 10091 19907
rect 10091 19873 10100 19907
rect 10048 19864 10100 19873
rect 11152 19907 11204 19916
rect 11152 19873 11161 19907
rect 11161 19873 11195 19907
rect 11195 19873 11204 19907
rect 11152 19864 11204 19873
rect 4252 19796 4304 19848
rect 4896 19796 4948 19848
rect 5172 19796 5224 19848
rect 9772 19839 9824 19848
rect 9772 19805 9781 19839
rect 9781 19805 9815 19839
rect 9815 19805 9824 19839
rect 9772 19796 9824 19805
rect 11612 19864 11664 19916
rect 5264 19728 5316 19780
rect 7104 19771 7156 19780
rect 7104 19737 7113 19771
rect 7113 19737 7147 19771
rect 7147 19737 7156 19771
rect 7104 19728 7156 19737
rect 12348 19839 12400 19848
rect 12348 19805 12357 19839
rect 12357 19805 12391 19839
rect 12391 19805 12400 19839
rect 12348 19796 12400 19805
rect 13360 19864 13412 19916
rect 14648 19864 14700 19916
rect 15752 19907 15804 19916
rect 15752 19873 15761 19907
rect 15761 19873 15795 19907
rect 15795 19873 15804 19907
rect 15752 19864 15804 19873
rect 18052 20000 18104 20052
rect 18236 20000 18288 20052
rect 18604 20000 18656 20052
rect 22008 20000 22060 20052
rect 15200 19796 15252 19848
rect 17224 19839 17276 19848
rect 17224 19805 17233 19839
rect 17233 19805 17267 19839
rect 17267 19805 17276 19839
rect 17224 19796 17276 19805
rect 18696 19975 18748 19984
rect 18696 19941 18705 19975
rect 18705 19941 18739 19975
rect 18739 19941 18748 19975
rect 18696 19932 18748 19941
rect 19984 19864 20036 19916
rect 20720 19864 20772 19916
rect 21272 19864 21324 19916
rect 21548 19864 21600 19916
rect 6920 19660 6972 19712
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 13820 19660 13872 19712
rect 18420 19703 18472 19712
rect 18420 19669 18429 19703
rect 18429 19669 18463 19703
rect 18463 19669 18472 19703
rect 18420 19660 18472 19669
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 19156 19703 19208 19712
rect 19156 19669 19165 19703
rect 19165 19669 19199 19703
rect 19199 19669 19208 19703
rect 19156 19660 19208 19669
rect 21088 19703 21140 19712
rect 21088 19669 21097 19703
rect 21097 19669 21131 19703
rect 21131 19669 21140 19703
rect 21088 19660 21140 19669
rect 22192 19660 22244 19712
rect 3662 19558 3714 19610
rect 3726 19558 3778 19610
rect 3790 19558 3842 19610
rect 3854 19558 3906 19610
rect 3918 19558 3970 19610
rect 5356 19456 5408 19508
rect 9128 19388 9180 19440
rect 4436 19252 4488 19304
rect 4896 19252 4948 19304
rect 8392 19320 8444 19372
rect 5724 19252 5776 19304
rect 5816 19295 5868 19304
rect 5816 19261 5825 19295
rect 5825 19261 5859 19295
rect 5859 19261 5868 19295
rect 5816 19252 5868 19261
rect 6000 19252 6052 19304
rect 7104 19295 7156 19304
rect 7104 19261 7113 19295
rect 7113 19261 7147 19295
rect 7147 19261 7156 19295
rect 7104 19252 7156 19261
rect 7288 19252 7340 19304
rect 8208 19252 8260 19304
rect 9772 19320 9824 19372
rect 10232 19295 10284 19304
rect 10232 19261 10241 19295
rect 10241 19261 10275 19295
rect 10275 19261 10284 19295
rect 10232 19252 10284 19261
rect 11152 19320 11204 19372
rect 12256 19456 12308 19508
rect 15752 19456 15804 19508
rect 12532 19388 12584 19440
rect 11520 19320 11572 19372
rect 11796 19363 11848 19372
rect 11796 19329 11805 19363
rect 11805 19329 11839 19363
rect 11839 19329 11848 19363
rect 11796 19320 11848 19329
rect 12164 19320 12216 19372
rect 13452 19320 13504 19372
rect 4712 19116 4764 19168
rect 4896 19116 4948 19168
rect 5356 19116 5408 19168
rect 5540 19159 5592 19168
rect 5540 19125 5549 19159
rect 5549 19125 5583 19159
rect 5583 19125 5592 19159
rect 5540 19116 5592 19125
rect 6920 19116 6972 19168
rect 10508 19184 10560 19236
rect 11428 19184 11480 19236
rect 14004 19320 14056 19372
rect 14096 19320 14148 19372
rect 17224 19388 17276 19440
rect 16672 19320 16724 19372
rect 15384 19295 15436 19304
rect 15384 19261 15393 19295
rect 15393 19261 15427 19295
rect 15427 19261 15436 19295
rect 15384 19252 15436 19261
rect 16304 19295 16356 19304
rect 16304 19261 16313 19295
rect 16313 19261 16347 19295
rect 16347 19261 16356 19295
rect 16304 19252 16356 19261
rect 18420 19320 18472 19372
rect 18880 19388 18932 19440
rect 19156 19388 19208 19440
rect 19984 19499 20036 19508
rect 19984 19465 19993 19499
rect 19993 19465 20027 19499
rect 20027 19465 20036 19499
rect 19984 19456 20036 19465
rect 21180 19456 21232 19508
rect 21456 19456 21508 19508
rect 21640 19456 21692 19508
rect 17684 19252 17736 19304
rect 18788 19184 18840 19236
rect 8392 19159 8444 19168
rect 8392 19125 8401 19159
rect 8401 19125 8435 19159
rect 8435 19125 8444 19159
rect 8392 19116 8444 19125
rect 12348 19116 12400 19168
rect 12716 19159 12768 19168
rect 12716 19125 12725 19159
rect 12725 19125 12759 19159
rect 12759 19125 12768 19159
rect 12716 19116 12768 19125
rect 17316 19116 17368 19168
rect 18052 19159 18104 19168
rect 18052 19125 18061 19159
rect 18061 19125 18095 19159
rect 18095 19125 18104 19159
rect 18052 19116 18104 19125
rect 18604 19116 18656 19168
rect 19524 19116 19576 19168
rect 20352 19295 20404 19304
rect 20352 19261 20361 19295
rect 20361 19261 20395 19295
rect 20395 19261 20404 19295
rect 20352 19252 20404 19261
rect 20628 19295 20680 19304
rect 20628 19261 20637 19295
rect 20637 19261 20671 19295
rect 20671 19261 20680 19295
rect 20628 19252 20680 19261
rect 20720 19252 20772 19304
rect 20812 19295 20864 19304
rect 20812 19261 20821 19295
rect 20821 19261 20855 19295
rect 20855 19261 20864 19295
rect 20812 19252 20864 19261
rect 21088 19320 21140 19372
rect 21364 19295 21416 19304
rect 21364 19261 21395 19295
rect 21395 19261 21416 19295
rect 21364 19252 21416 19261
rect 22284 19295 22336 19304
rect 22284 19261 22293 19295
rect 22293 19261 22327 19295
rect 22327 19261 22336 19295
rect 22284 19252 22336 19261
rect 22192 19227 22244 19236
rect 22192 19193 22201 19227
rect 22201 19193 22235 19227
rect 22235 19193 22244 19227
rect 22192 19184 22244 19193
rect 20444 19116 20496 19168
rect 20720 19116 20772 19168
rect 20996 19116 21048 19168
rect 21824 19159 21876 19168
rect 21824 19125 21833 19159
rect 21833 19125 21867 19159
rect 21867 19125 21876 19159
rect 21824 19116 21876 19125
rect 22100 19116 22152 19168
rect 19022 19014 19074 19066
rect 19086 19014 19138 19066
rect 19150 19014 19202 19066
rect 19214 19014 19266 19066
rect 19278 19014 19330 19066
rect 5540 18912 5592 18964
rect 5724 18912 5776 18964
rect 7932 18912 7984 18964
rect 8392 18912 8444 18964
rect 4712 18776 4764 18828
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 6828 18819 6880 18828
rect 6828 18785 6837 18819
rect 6837 18785 6871 18819
rect 6871 18785 6880 18819
rect 6828 18776 6880 18785
rect 8300 18844 8352 18896
rect 8208 18819 8260 18828
rect 8208 18785 8217 18819
rect 8217 18785 8251 18819
rect 8251 18785 8260 18819
rect 8208 18776 8260 18785
rect 8760 18776 8812 18828
rect 10048 18912 10100 18964
rect 10876 18912 10928 18964
rect 9128 18844 9180 18896
rect 9404 18776 9456 18828
rect 6000 18708 6052 18760
rect 9864 18708 9916 18760
rect 10508 18776 10560 18828
rect 15200 18912 15252 18964
rect 18052 18912 18104 18964
rect 18604 18912 18656 18964
rect 17684 18844 17736 18896
rect 11796 18640 11848 18692
rect 12256 18708 12308 18760
rect 14740 18776 14792 18828
rect 14924 18776 14976 18828
rect 16488 18776 16540 18828
rect 19156 18912 19208 18964
rect 19294 18912 19346 18964
rect 20352 18912 20404 18964
rect 21180 18912 21232 18964
rect 22560 18912 22612 18964
rect 18788 18776 18840 18828
rect 19156 18819 19208 18828
rect 19156 18785 19197 18819
rect 19197 18785 19208 18819
rect 19156 18776 19208 18785
rect 19294 18776 19346 18828
rect 21364 18819 21416 18828
rect 21364 18785 21373 18819
rect 21373 18785 21407 18819
rect 21407 18785 21416 18819
rect 21364 18776 21416 18785
rect 22192 18819 22244 18828
rect 22192 18785 22201 18819
rect 22201 18785 22235 18819
rect 22235 18785 22244 18819
rect 22192 18776 22244 18785
rect 16396 18708 16448 18760
rect 17316 18708 17368 18760
rect 12440 18640 12492 18692
rect 6460 18615 6512 18624
rect 6460 18581 6469 18615
rect 6469 18581 6503 18615
rect 6503 18581 6512 18615
rect 6460 18572 6512 18581
rect 7840 18572 7892 18624
rect 9496 18615 9548 18624
rect 9496 18581 9505 18615
rect 9505 18581 9539 18615
rect 9539 18581 9548 18615
rect 9496 18572 9548 18581
rect 12256 18615 12308 18624
rect 12256 18581 12265 18615
rect 12265 18581 12299 18615
rect 12299 18581 12308 18615
rect 12256 18572 12308 18581
rect 12348 18572 12400 18624
rect 13084 18572 13136 18624
rect 18696 18640 18748 18692
rect 18788 18615 18840 18624
rect 18788 18581 18797 18615
rect 18797 18581 18831 18615
rect 18831 18581 18840 18615
rect 18788 18572 18840 18581
rect 18972 18572 19024 18624
rect 19156 18572 19208 18624
rect 19432 18708 19484 18760
rect 20628 18708 20680 18760
rect 21088 18708 21140 18760
rect 20444 18615 20496 18624
rect 20444 18581 20453 18615
rect 20453 18581 20487 18615
rect 20487 18581 20496 18615
rect 20444 18572 20496 18581
rect 20628 18615 20680 18624
rect 20628 18581 20637 18615
rect 20637 18581 20671 18615
rect 20671 18581 20680 18615
rect 20628 18572 20680 18581
rect 21364 18572 21416 18624
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 6092 18368 6144 18420
rect 6920 18368 6972 18420
rect 4252 18164 4304 18216
rect 5264 18232 5316 18284
rect 5356 18232 5408 18284
rect 6000 18275 6052 18284
rect 6000 18241 6009 18275
rect 6009 18241 6043 18275
rect 6043 18241 6052 18275
rect 6000 18232 6052 18241
rect 5724 18164 5776 18216
rect 5816 18139 5868 18148
rect 5816 18105 5825 18139
rect 5825 18105 5859 18139
rect 5859 18105 5868 18139
rect 6460 18164 6512 18216
rect 6920 18232 6972 18284
rect 8760 18368 8812 18420
rect 11796 18411 11848 18420
rect 11796 18377 11805 18411
rect 11805 18377 11839 18411
rect 11839 18377 11848 18411
rect 11796 18368 11848 18377
rect 14740 18368 14792 18420
rect 8208 18232 8260 18284
rect 9128 18232 9180 18284
rect 9404 18164 9456 18216
rect 10876 18275 10928 18284
rect 10876 18241 10885 18275
rect 10885 18241 10919 18275
rect 10919 18241 10928 18275
rect 10876 18232 10928 18241
rect 5816 18096 5868 18105
rect 8300 18096 8352 18148
rect 10968 18096 11020 18148
rect 12256 18232 12308 18284
rect 13084 18300 13136 18352
rect 12716 18232 12768 18284
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 12440 18164 12492 18216
rect 13544 18207 13596 18216
rect 13544 18173 13553 18207
rect 13553 18173 13587 18207
rect 13587 18173 13596 18207
rect 13544 18164 13596 18173
rect 13728 18207 13780 18216
rect 13728 18173 13737 18207
rect 13737 18173 13771 18207
rect 13771 18173 13780 18207
rect 13728 18164 13780 18173
rect 13912 18164 13964 18216
rect 12348 18096 12400 18148
rect 14924 18368 14976 18420
rect 20444 18368 20496 18420
rect 15936 18164 15988 18216
rect 16488 18300 16540 18352
rect 16396 18164 16448 18216
rect 21640 18368 21692 18420
rect 21824 18368 21876 18420
rect 22100 18368 22152 18420
rect 20720 18300 20772 18352
rect 22652 18300 22704 18352
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 17316 18207 17368 18216
rect 17316 18173 17325 18207
rect 17325 18173 17359 18207
rect 17359 18173 17368 18207
rect 17316 18164 17368 18173
rect 20720 18207 20772 18216
rect 20720 18173 20729 18207
rect 20729 18173 20763 18207
rect 20763 18173 20772 18207
rect 20720 18164 20772 18173
rect 20812 18207 20864 18216
rect 20812 18173 20821 18207
rect 20821 18173 20855 18207
rect 20855 18173 20864 18207
rect 20812 18164 20864 18173
rect 21456 18207 21508 18216
rect 21456 18173 21468 18207
rect 21468 18173 21502 18207
rect 21502 18173 21508 18207
rect 21456 18164 21508 18173
rect 4896 18028 4948 18080
rect 7380 18071 7432 18080
rect 7380 18037 7389 18071
rect 7389 18037 7423 18071
rect 7423 18037 7432 18071
rect 7380 18028 7432 18037
rect 8392 18071 8444 18080
rect 8392 18037 8401 18071
rect 8401 18037 8435 18071
rect 8435 18037 8444 18071
rect 8392 18028 8444 18037
rect 14556 18028 14608 18080
rect 16856 18096 16908 18148
rect 21364 18096 21416 18148
rect 16580 18028 16632 18080
rect 20352 18071 20404 18080
rect 20352 18037 20361 18071
rect 20361 18037 20395 18071
rect 20395 18037 20404 18071
rect 20352 18028 20404 18037
rect 21824 18096 21876 18148
rect 21640 18071 21692 18080
rect 21640 18037 21649 18071
rect 21649 18037 21683 18071
rect 21683 18037 21692 18071
rect 21640 18028 21692 18037
rect 21732 18028 21784 18080
rect 19022 17926 19074 17978
rect 19086 17926 19138 17978
rect 19150 17926 19202 17978
rect 19214 17926 19266 17978
rect 19278 17926 19330 17978
rect 6000 17824 6052 17876
rect 8300 17867 8352 17876
rect 8300 17833 8309 17867
rect 8309 17833 8343 17867
rect 8343 17833 8352 17867
rect 8300 17824 8352 17833
rect 4896 17688 4948 17740
rect 5816 17688 5868 17740
rect 6460 17688 6512 17740
rect 7380 17688 7432 17740
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 8208 17731 8260 17740
rect 8208 17697 8217 17731
rect 8217 17697 8251 17731
rect 8251 17697 8260 17731
rect 8208 17688 8260 17697
rect 13728 17824 13780 17876
rect 13820 17824 13872 17876
rect 15936 17824 15988 17876
rect 18788 17824 18840 17876
rect 19616 17867 19668 17876
rect 19616 17833 19631 17867
rect 19631 17833 19665 17867
rect 19665 17833 19668 17867
rect 19616 17824 19668 17833
rect 20812 17824 20864 17876
rect 21456 17824 21508 17876
rect 21824 17824 21876 17876
rect 9404 17688 9456 17740
rect 9864 17688 9916 17740
rect 10876 17688 10928 17740
rect 11244 17688 11296 17740
rect 13544 17731 13596 17740
rect 13544 17697 13550 17731
rect 13550 17697 13584 17731
rect 13584 17697 13596 17731
rect 13544 17688 13596 17697
rect 13912 17620 13964 17672
rect 14096 17620 14148 17672
rect 19340 17756 19392 17808
rect 19432 17756 19484 17808
rect 16396 17663 16448 17672
rect 16396 17629 16405 17663
rect 16405 17629 16439 17663
rect 16439 17629 16448 17663
rect 16396 17620 16448 17629
rect 19064 17731 19116 17740
rect 19064 17697 19073 17731
rect 19073 17697 19107 17731
rect 19107 17697 19116 17731
rect 19064 17688 19116 17697
rect 19156 17731 19208 17740
rect 19156 17697 19165 17731
rect 19165 17697 19199 17731
rect 19199 17697 19208 17731
rect 19156 17688 19208 17697
rect 15108 17552 15160 17604
rect 18972 17552 19024 17604
rect 20260 17731 20312 17740
rect 20260 17697 20269 17731
rect 20269 17697 20303 17731
rect 20303 17697 20312 17731
rect 20260 17688 20312 17697
rect 20996 17688 21048 17740
rect 21732 17756 21784 17808
rect 22284 17756 22336 17808
rect 21364 17688 21416 17740
rect 21548 17688 21600 17740
rect 20536 17620 20588 17672
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 23020 17663 23072 17672
rect 23020 17629 23029 17663
rect 23029 17629 23063 17663
rect 23063 17629 23072 17663
rect 23020 17620 23072 17629
rect 21364 17552 21416 17604
rect 7748 17527 7800 17536
rect 7748 17493 7757 17527
rect 7757 17493 7791 17527
rect 7791 17493 7800 17527
rect 7748 17484 7800 17493
rect 10048 17484 10100 17536
rect 11520 17527 11572 17536
rect 11520 17493 11529 17527
rect 11529 17493 11563 17527
rect 11563 17493 11572 17527
rect 11520 17484 11572 17493
rect 11980 17527 12032 17536
rect 11980 17493 11989 17527
rect 11989 17493 12023 17527
rect 12023 17493 12032 17527
rect 11980 17484 12032 17493
rect 14280 17484 14332 17536
rect 16212 17527 16264 17536
rect 16212 17493 16221 17527
rect 16221 17493 16255 17527
rect 16255 17493 16264 17527
rect 16212 17484 16264 17493
rect 18236 17484 18288 17536
rect 19156 17484 19208 17536
rect 20628 17484 20680 17536
rect 21088 17527 21140 17536
rect 21088 17493 21097 17527
rect 21097 17493 21131 17527
rect 21131 17493 21140 17527
rect 21088 17484 21140 17493
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 7748 17280 7800 17332
rect 11980 17280 12032 17332
rect 12164 17280 12216 17332
rect 14280 17280 14332 17332
rect 16212 17280 16264 17332
rect 16672 17280 16724 17332
rect 18788 17280 18840 17332
rect 18972 17280 19024 17332
rect 19064 17280 19116 17332
rect 21088 17280 21140 17332
rect 21364 17280 21416 17332
rect 8208 17144 8260 17196
rect 9404 17076 9456 17128
rect 10048 17144 10100 17196
rect 11520 17144 11572 17196
rect 14280 17144 14332 17196
rect 11152 17008 11204 17060
rect 13820 17076 13872 17128
rect 14096 17076 14148 17128
rect 14556 17076 14608 17128
rect 14740 17187 14792 17196
rect 14740 17153 14749 17187
rect 14749 17153 14783 17187
rect 14783 17153 14792 17187
rect 14740 17144 14792 17153
rect 17500 17212 17552 17264
rect 12532 17008 12584 17060
rect 13176 17008 13228 17060
rect 13268 17008 13320 17060
rect 14188 17008 14240 17060
rect 15936 17008 15988 17060
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 16948 17051 17000 17060
rect 16948 17017 16957 17051
rect 16957 17017 16991 17051
rect 16991 17017 17000 17051
rect 16948 17008 17000 17017
rect 9220 16983 9272 16992
rect 9220 16949 9229 16983
rect 9229 16949 9263 16983
rect 9263 16949 9272 16983
rect 9220 16940 9272 16949
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 11428 16940 11480 16992
rect 11704 16983 11756 16992
rect 11704 16949 11713 16983
rect 11713 16949 11747 16983
rect 11747 16949 11756 16983
rect 11704 16940 11756 16949
rect 12164 16940 12216 16992
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 15016 16940 15068 16992
rect 16764 16940 16816 16992
rect 17132 16940 17184 16992
rect 18236 17008 18288 17060
rect 22192 17212 22244 17264
rect 19800 17076 19852 17128
rect 20352 17076 20404 17128
rect 20536 17076 20588 17128
rect 21180 17119 21232 17128
rect 21180 17085 21189 17119
rect 21189 17085 21223 17119
rect 21223 17085 21232 17119
rect 21180 17076 21232 17085
rect 21732 17076 21784 17128
rect 20076 16940 20128 16992
rect 19022 16838 19074 16890
rect 19086 16838 19138 16890
rect 19150 16838 19202 16890
rect 19214 16838 19266 16890
rect 19278 16838 19330 16890
rect 7012 16736 7064 16788
rect 6460 16600 6512 16652
rect 6184 16532 6236 16584
rect 6828 16600 6880 16652
rect 9220 16668 9272 16720
rect 10784 16736 10836 16788
rect 11520 16779 11572 16788
rect 11520 16745 11529 16779
rect 11529 16745 11563 16779
rect 11563 16745 11572 16779
rect 11520 16736 11572 16745
rect 12532 16779 12584 16788
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 13268 16736 13320 16788
rect 14740 16779 14792 16788
rect 14740 16745 14749 16779
rect 14749 16745 14783 16779
rect 14783 16745 14792 16779
rect 14740 16736 14792 16745
rect 16856 16736 16908 16788
rect 17408 16736 17460 16788
rect 19432 16736 19484 16788
rect 22652 16779 22704 16788
rect 22652 16745 22661 16779
rect 22661 16745 22695 16779
rect 22695 16745 22704 16779
rect 22652 16736 22704 16745
rect 11060 16600 11112 16652
rect 11152 16600 11204 16652
rect 11428 16600 11480 16652
rect 12624 16643 12676 16652
rect 12624 16609 12634 16643
rect 12634 16609 12676 16643
rect 12624 16600 12676 16609
rect 11888 16532 11940 16584
rect 13084 16532 13136 16584
rect 13176 16532 13228 16584
rect 9496 16464 9548 16516
rect 6552 16396 6604 16448
rect 6644 16439 6696 16448
rect 6644 16405 6653 16439
rect 6653 16405 6687 16439
rect 6687 16405 6696 16439
rect 6644 16396 6696 16405
rect 6920 16396 6972 16448
rect 15660 16600 15712 16652
rect 16580 16600 16632 16652
rect 17132 16600 17184 16652
rect 21640 16668 21692 16720
rect 14372 16532 14424 16584
rect 12164 16439 12216 16448
rect 12164 16405 12173 16439
rect 12173 16405 12207 16439
rect 12207 16405 12216 16439
rect 12164 16396 12216 16405
rect 13912 16396 13964 16448
rect 14648 16439 14700 16448
rect 14648 16405 14657 16439
rect 14657 16405 14691 16439
rect 14691 16405 14700 16439
rect 14648 16396 14700 16405
rect 14924 16396 14976 16448
rect 16856 16532 16908 16584
rect 17040 16575 17092 16584
rect 17040 16541 17049 16575
rect 17049 16541 17083 16575
rect 17083 16541 17092 16575
rect 19616 16600 19668 16652
rect 19800 16600 19852 16652
rect 23020 16600 23072 16652
rect 17040 16532 17092 16541
rect 16672 16464 16724 16516
rect 21180 16532 21232 16584
rect 16580 16396 16632 16448
rect 16948 16396 17000 16448
rect 18880 16396 18932 16448
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 6184 16192 6236 16244
rect 9496 16192 9548 16244
rect 6460 16124 6512 16176
rect 5080 16031 5132 16040
rect 5080 15997 5089 16031
rect 5089 15997 5123 16031
rect 5123 15997 5132 16031
rect 6368 16056 6420 16108
rect 6920 16056 6972 16108
rect 5080 15988 5132 15997
rect 5540 15963 5592 15972
rect 5540 15929 5549 15963
rect 5549 15929 5583 15963
rect 5583 15929 5592 15963
rect 5540 15920 5592 15929
rect 5908 15988 5960 16040
rect 6460 16031 6512 16040
rect 6460 15997 6469 16031
rect 6469 15997 6503 16031
rect 6503 15997 6512 16031
rect 6460 15988 6512 15997
rect 6644 15988 6696 16040
rect 6092 15963 6144 15972
rect 6092 15929 6101 15963
rect 6101 15929 6135 15963
rect 6135 15929 6144 15963
rect 6092 15920 6144 15929
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 5448 15852 5500 15904
rect 5632 15852 5684 15904
rect 6000 15852 6052 15904
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 8024 16056 8076 16108
rect 11152 16099 11204 16108
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 11152 16056 11204 16065
rect 7840 15988 7892 16040
rect 9220 15988 9272 16040
rect 11428 15988 11480 16040
rect 13912 16031 13964 16040
rect 13912 15997 13921 16031
rect 13921 15997 13955 16031
rect 13955 15997 13964 16031
rect 13912 15988 13964 15997
rect 15108 16192 15160 16244
rect 22100 16192 22152 16244
rect 14648 16124 14700 16176
rect 14372 16031 14424 16040
rect 14372 15997 14381 16031
rect 14381 15997 14415 16031
rect 14415 15997 14424 16031
rect 14372 15988 14424 15997
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 16580 16124 16632 16176
rect 23020 16192 23072 16244
rect 15016 16099 15068 16108
rect 15016 16065 15025 16099
rect 15025 16065 15059 16099
rect 15059 16065 15068 16099
rect 15016 16056 15068 16065
rect 15108 16031 15160 16040
rect 15108 15997 15117 16031
rect 15117 15997 15151 16031
rect 15151 15997 15160 16031
rect 15108 15988 15160 15997
rect 15936 15988 15988 16040
rect 16396 15988 16448 16040
rect 16672 15988 16724 16040
rect 16764 16031 16816 16040
rect 16764 15997 16773 16031
rect 16773 15997 16807 16031
rect 16807 15997 16816 16031
rect 16764 15988 16816 15997
rect 17040 16031 17092 16040
rect 17040 15997 17049 16031
rect 17049 15997 17083 16031
rect 17083 15997 17092 16031
rect 17040 15988 17092 15997
rect 22376 16056 22428 16108
rect 22836 15988 22888 16040
rect 6736 15852 6788 15904
rect 7288 15852 7340 15904
rect 7656 15852 7708 15904
rect 9864 15895 9916 15904
rect 9864 15861 9873 15895
rect 9873 15861 9907 15895
rect 9907 15861 9916 15895
rect 9864 15852 9916 15861
rect 10416 15895 10468 15904
rect 10416 15861 10425 15895
rect 10425 15861 10459 15895
rect 10459 15861 10468 15895
rect 10416 15852 10468 15861
rect 11796 15895 11848 15904
rect 11796 15861 11805 15895
rect 11805 15861 11839 15895
rect 11839 15861 11848 15895
rect 11796 15852 11848 15861
rect 18236 15920 18288 15972
rect 22008 15920 22060 15972
rect 15476 15895 15528 15904
rect 15476 15861 15485 15895
rect 15485 15861 15519 15895
rect 15519 15861 15528 15895
rect 15476 15852 15528 15861
rect 15660 15895 15712 15904
rect 15660 15861 15669 15895
rect 15669 15861 15703 15895
rect 15703 15861 15712 15895
rect 15660 15852 15712 15861
rect 17408 15895 17460 15904
rect 17408 15861 17417 15895
rect 17417 15861 17451 15895
rect 17451 15861 17460 15895
rect 17408 15852 17460 15861
rect 19022 15750 19074 15802
rect 19086 15750 19138 15802
rect 19150 15750 19202 15802
rect 19214 15750 19266 15802
rect 19278 15750 19330 15802
rect 5172 15648 5224 15700
rect 5540 15648 5592 15700
rect 5908 15648 5960 15700
rect 6092 15648 6144 15700
rect 9864 15648 9916 15700
rect 10416 15648 10468 15700
rect 6552 15580 6604 15632
rect 5540 15512 5592 15564
rect 6184 15555 6236 15564
rect 6184 15521 6193 15555
rect 6193 15521 6227 15555
rect 6227 15521 6236 15555
rect 6184 15512 6236 15521
rect 6368 15512 6420 15564
rect 6736 15555 6788 15564
rect 6736 15521 6745 15555
rect 6745 15521 6779 15555
rect 6779 15521 6788 15555
rect 6736 15512 6788 15521
rect 6828 15512 6880 15564
rect 7288 15580 7340 15632
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 7840 15487 7892 15496
rect 7840 15453 7849 15487
rect 7849 15453 7883 15487
rect 7883 15453 7892 15487
rect 7840 15444 7892 15453
rect 8024 15555 8076 15564
rect 8024 15521 8033 15555
rect 8033 15521 8067 15555
rect 8067 15521 8076 15555
rect 8024 15512 8076 15521
rect 14372 15648 14424 15700
rect 16396 15648 16448 15700
rect 18880 15648 18932 15700
rect 20076 15691 20128 15700
rect 20076 15657 20085 15691
rect 20085 15657 20119 15691
rect 20119 15657 20128 15691
rect 20076 15648 20128 15657
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 11060 15487 11112 15496
rect 11060 15453 11069 15487
rect 11069 15453 11103 15487
rect 11103 15453 11112 15487
rect 11060 15444 11112 15453
rect 12992 15512 13044 15564
rect 13176 15555 13228 15564
rect 13176 15521 13185 15555
rect 13185 15521 13219 15555
rect 13219 15521 13228 15555
rect 13176 15512 13228 15521
rect 13452 15555 13504 15564
rect 13452 15521 13461 15555
rect 13461 15521 13495 15555
rect 13495 15521 13504 15555
rect 13452 15512 13504 15521
rect 12532 15444 12584 15496
rect 4528 15308 4580 15360
rect 6000 15308 6052 15360
rect 7196 15351 7248 15360
rect 7196 15317 7205 15351
rect 7205 15317 7239 15351
rect 7239 15317 7248 15351
rect 7196 15308 7248 15317
rect 7748 15308 7800 15360
rect 8208 15351 8260 15360
rect 8208 15317 8217 15351
rect 8217 15317 8251 15351
rect 8251 15317 8260 15351
rect 8208 15308 8260 15317
rect 8300 15351 8352 15360
rect 8300 15317 8309 15351
rect 8309 15317 8343 15351
rect 8343 15317 8352 15351
rect 8300 15308 8352 15317
rect 14556 15512 14608 15564
rect 14648 15512 14700 15564
rect 14924 15512 14976 15564
rect 21180 15580 21232 15632
rect 22836 15580 22888 15632
rect 16672 15512 16724 15564
rect 18420 15512 18472 15564
rect 19984 15555 20036 15564
rect 19984 15521 19993 15555
rect 19993 15521 20027 15555
rect 20027 15521 20036 15555
rect 19984 15512 20036 15521
rect 15660 15444 15712 15496
rect 15200 15419 15252 15428
rect 15200 15385 15209 15419
rect 15209 15385 15243 15419
rect 15243 15385 15252 15419
rect 15200 15376 15252 15385
rect 17040 15487 17092 15496
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 17776 15444 17828 15496
rect 19432 15444 19484 15496
rect 21364 15512 21416 15564
rect 9036 15308 9088 15360
rect 9864 15351 9916 15360
rect 9864 15317 9873 15351
rect 9873 15317 9907 15351
rect 9907 15317 9916 15351
rect 9864 15308 9916 15317
rect 11428 15351 11480 15360
rect 11428 15317 11437 15351
rect 11437 15317 11471 15351
rect 11471 15317 11480 15351
rect 11428 15308 11480 15317
rect 16580 15308 16632 15360
rect 19524 15351 19576 15360
rect 19524 15317 19533 15351
rect 19533 15317 19567 15351
rect 19567 15317 19576 15351
rect 19524 15308 19576 15317
rect 19616 15351 19668 15360
rect 19616 15317 19625 15351
rect 19625 15317 19659 15351
rect 19659 15317 19668 15351
rect 19616 15308 19668 15317
rect 22008 15308 22060 15360
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 6460 15104 6512 15156
rect 6920 15104 6972 15156
rect 7196 15104 7248 15156
rect 8300 15104 8352 15156
rect 11428 15104 11480 15156
rect 13452 15104 13504 15156
rect 17776 15147 17828 15156
rect 17776 15113 17785 15147
rect 17785 15113 17819 15147
rect 17819 15113 17828 15147
rect 17776 15104 17828 15113
rect 7748 15036 7800 15088
rect 6644 15011 6696 15020
rect 6644 14977 6653 15011
rect 6653 14977 6687 15011
rect 6687 14977 6696 15011
rect 6644 14968 6696 14977
rect 4528 14900 4580 14952
rect 5632 14900 5684 14952
rect 6920 14943 6972 14952
rect 6920 14909 6929 14943
rect 6929 14909 6963 14943
rect 6963 14909 6972 14943
rect 6920 14900 6972 14909
rect 8392 14968 8444 15020
rect 8208 14943 8260 14952
rect 8208 14909 8217 14943
rect 8217 14909 8251 14943
rect 8251 14909 8260 14943
rect 8208 14900 8260 14909
rect 9036 14943 9088 14952
rect 9036 14909 9045 14943
rect 9045 14909 9079 14943
rect 9079 14909 9088 14943
rect 9036 14900 9088 14909
rect 12164 15036 12216 15088
rect 13912 15036 13964 15088
rect 11704 14968 11756 15020
rect 12072 14968 12124 15020
rect 11520 14943 11572 14952
rect 11520 14909 11529 14943
rect 11529 14909 11563 14943
rect 11563 14909 11572 14943
rect 11520 14900 11572 14909
rect 11796 14900 11848 14952
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 8300 14832 8352 14884
rect 12808 14875 12860 14884
rect 12808 14841 12817 14875
rect 12817 14841 12851 14875
rect 12851 14841 12860 14875
rect 12808 14832 12860 14841
rect 13084 14832 13136 14884
rect 6736 14764 6788 14816
rect 7012 14807 7064 14816
rect 7012 14773 7021 14807
rect 7021 14773 7055 14807
rect 7055 14773 7064 14807
rect 7012 14764 7064 14773
rect 7104 14764 7156 14816
rect 7840 14764 7892 14816
rect 8116 14764 8168 14816
rect 9128 14807 9180 14816
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 11888 14807 11940 14816
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 11980 14764 12032 14816
rect 12348 14764 12400 14816
rect 14188 14943 14240 14952
rect 14188 14909 14197 14943
rect 14197 14909 14231 14943
rect 14231 14909 14240 14943
rect 14188 14900 14240 14909
rect 16396 14900 16448 14952
rect 16580 14943 16632 14952
rect 16580 14909 16614 14943
rect 16614 14909 16632 14943
rect 16580 14900 16632 14909
rect 13728 14764 13780 14816
rect 17684 14807 17736 14816
rect 17684 14773 17693 14807
rect 17693 14773 17727 14807
rect 17727 14773 17736 14807
rect 19616 15104 19668 15156
rect 19984 15104 20036 15156
rect 21364 15147 21416 15156
rect 21364 15113 21373 15147
rect 21373 15113 21407 15147
rect 21407 15113 21416 15147
rect 21364 15104 21416 15113
rect 18696 14943 18748 14952
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 19524 14900 19576 14952
rect 20720 14900 20772 14952
rect 21916 15011 21968 15020
rect 21916 14977 21925 15011
rect 21925 14977 21959 15011
rect 21959 14977 21968 15011
rect 21916 14968 21968 14977
rect 22008 14900 22060 14952
rect 20260 14832 20312 14884
rect 22652 14900 22704 14952
rect 22468 14875 22520 14884
rect 22468 14841 22477 14875
rect 22477 14841 22511 14875
rect 22511 14841 22520 14875
rect 22468 14832 22520 14841
rect 17684 14764 17736 14773
rect 19524 14764 19576 14816
rect 20168 14807 20220 14816
rect 20168 14773 20177 14807
rect 20177 14773 20211 14807
rect 20211 14773 20220 14807
rect 20168 14764 20220 14773
rect 21456 14764 21508 14816
rect 22376 14764 22428 14816
rect 19022 14662 19074 14714
rect 19086 14662 19138 14714
rect 19150 14662 19202 14714
rect 19214 14662 19266 14714
rect 19278 14662 19330 14714
rect 4896 14560 4948 14612
rect 5724 14424 5776 14476
rect 6736 14560 6788 14612
rect 7012 14560 7064 14612
rect 9404 14560 9456 14612
rect 7840 14492 7892 14544
rect 11980 14560 12032 14612
rect 12072 14560 12124 14612
rect 6644 14467 6696 14476
rect 6644 14433 6653 14467
rect 6653 14433 6687 14467
rect 6687 14433 6696 14467
rect 6644 14424 6696 14433
rect 6736 14467 6788 14476
rect 6736 14433 6745 14467
rect 6745 14433 6779 14467
rect 6779 14433 6788 14467
rect 6736 14424 6788 14433
rect 7104 14424 7156 14476
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 7380 14473 7432 14482
rect 7380 14439 7389 14473
rect 7389 14439 7423 14473
rect 7423 14439 7432 14473
rect 7380 14430 7432 14439
rect 7472 14470 7524 14476
rect 7472 14436 7484 14470
rect 7484 14436 7518 14470
rect 7518 14436 7524 14470
rect 7472 14424 7524 14436
rect 7748 14424 7800 14476
rect 9864 14467 9916 14476
rect 9864 14433 9876 14467
rect 9876 14433 9910 14467
rect 9910 14433 9916 14467
rect 9864 14424 9916 14433
rect 5448 14356 5500 14408
rect 7288 14356 7340 14408
rect 8300 14356 8352 14408
rect 9128 14356 9180 14408
rect 4252 14220 4304 14272
rect 6644 14288 6696 14340
rect 8116 14331 8168 14340
rect 8116 14297 8125 14331
rect 8125 14297 8159 14331
rect 8159 14297 8168 14331
rect 8116 14288 8168 14297
rect 9496 14331 9548 14340
rect 9496 14297 9505 14331
rect 9505 14297 9539 14331
rect 9539 14297 9548 14331
rect 11704 14424 11756 14476
rect 12808 14560 12860 14612
rect 13176 14560 13228 14612
rect 13912 14560 13964 14612
rect 14188 14560 14240 14612
rect 17408 14560 17460 14612
rect 18420 14603 18472 14612
rect 18420 14569 18429 14603
rect 18429 14569 18463 14603
rect 18463 14569 18472 14603
rect 18420 14560 18472 14569
rect 20168 14560 20220 14612
rect 12532 14492 12584 14544
rect 13084 14492 13136 14544
rect 12440 14467 12492 14476
rect 12440 14433 12449 14467
rect 12449 14433 12483 14467
rect 12483 14433 12492 14467
rect 12440 14424 12492 14433
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 11612 14356 11664 14408
rect 9496 14288 9548 14297
rect 10968 14331 11020 14340
rect 10968 14297 10977 14331
rect 10977 14297 11011 14331
rect 11011 14297 11020 14331
rect 16396 14492 16448 14544
rect 21640 14560 21692 14612
rect 22468 14560 22520 14612
rect 17776 14424 17828 14476
rect 18696 14424 18748 14476
rect 19708 14424 19760 14476
rect 15844 14356 15896 14408
rect 21456 14467 21508 14476
rect 21456 14433 21465 14467
rect 21465 14433 21499 14467
rect 21499 14433 21508 14467
rect 21456 14424 21508 14433
rect 10968 14288 11020 14297
rect 13268 14288 13320 14340
rect 7196 14220 7248 14272
rect 7840 14263 7892 14272
rect 7840 14229 7849 14263
rect 7849 14229 7883 14263
rect 7883 14229 7892 14263
rect 7840 14220 7892 14229
rect 7932 14263 7984 14272
rect 7932 14229 7941 14263
rect 7941 14229 7975 14263
rect 7975 14229 7984 14263
rect 7932 14220 7984 14229
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 11888 14220 11940 14272
rect 13728 14220 13780 14272
rect 13820 14263 13872 14272
rect 13820 14229 13829 14263
rect 13829 14229 13863 14263
rect 13863 14229 13872 14263
rect 13820 14220 13872 14229
rect 16764 14220 16816 14272
rect 20996 14356 21048 14408
rect 21548 14399 21600 14408
rect 21548 14365 21557 14399
rect 21557 14365 21591 14399
rect 21591 14365 21600 14399
rect 21548 14356 21600 14365
rect 22100 14467 22152 14476
rect 22100 14433 22109 14467
rect 22109 14433 22143 14467
rect 22143 14433 22152 14467
rect 22100 14424 22152 14433
rect 21456 14288 21508 14340
rect 19432 14220 19484 14272
rect 21180 14220 21232 14272
rect 22192 14220 22244 14272
rect 22468 14263 22520 14272
rect 22468 14229 22477 14263
rect 22477 14229 22511 14263
rect 22511 14229 22520 14263
rect 22468 14220 22520 14229
rect 22652 14220 22704 14272
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 5724 14059 5776 14068
rect 5724 14025 5733 14059
rect 5733 14025 5767 14059
rect 5767 14025 5776 14059
rect 5724 14016 5776 14025
rect 7196 14016 7248 14068
rect 9864 14016 9916 14068
rect 11428 14016 11480 14068
rect 12440 14016 12492 14068
rect 13820 14016 13872 14068
rect 10232 13948 10284 14000
rect 7932 13880 7984 13932
rect 8208 13880 8260 13932
rect 11428 13923 11480 13932
rect 11428 13889 11437 13923
rect 11437 13889 11471 13923
rect 11471 13889 11480 13923
rect 11428 13880 11480 13889
rect 13268 13880 13320 13932
rect 15200 13880 15252 13932
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 16396 13880 16448 13932
rect 4436 13812 4488 13864
rect 6736 13812 6788 13864
rect 8300 13812 8352 13864
rect 4160 13744 4212 13796
rect 9404 13855 9456 13864
rect 9404 13821 9413 13855
rect 9413 13821 9447 13855
rect 9447 13821 9456 13855
rect 9404 13812 9456 13821
rect 11704 13812 11756 13864
rect 13084 13812 13136 13864
rect 10048 13744 10100 13796
rect 10968 13744 11020 13796
rect 13728 13855 13780 13864
rect 13728 13821 13737 13855
rect 13737 13821 13771 13855
rect 13771 13821 13780 13855
rect 13728 13812 13780 13821
rect 16028 13855 16080 13864
rect 16028 13821 16037 13855
rect 16037 13821 16071 13855
rect 16071 13821 16080 13855
rect 16028 13812 16080 13821
rect 16120 13744 16172 13796
rect 16764 14016 16816 14068
rect 17040 14016 17092 14068
rect 17776 14016 17828 14068
rect 19432 14016 19484 14068
rect 21456 14016 21508 14068
rect 22192 14016 22244 14068
rect 20720 13948 20772 14000
rect 21180 13923 21232 13932
rect 21180 13889 21189 13923
rect 21189 13889 21223 13923
rect 21223 13889 21232 13923
rect 21180 13880 21232 13889
rect 21456 13923 21508 13932
rect 21456 13889 21465 13923
rect 21465 13889 21499 13923
rect 21499 13889 21508 13923
rect 21456 13880 21508 13889
rect 19340 13812 19392 13864
rect 19524 13812 19576 13864
rect 20352 13812 20404 13864
rect 20536 13812 20588 13864
rect 20996 13812 21048 13864
rect 22100 13812 22152 13864
rect 20444 13787 20496 13796
rect 20444 13753 20453 13787
rect 20453 13753 20487 13787
rect 20487 13753 20496 13787
rect 20444 13744 20496 13753
rect 8576 13676 8628 13728
rect 9772 13719 9824 13728
rect 9772 13685 9781 13719
rect 9781 13685 9815 13719
rect 9815 13685 9824 13719
rect 9772 13676 9824 13685
rect 11796 13719 11848 13728
rect 11796 13685 11805 13719
rect 11805 13685 11839 13719
rect 11839 13685 11848 13719
rect 11796 13676 11848 13685
rect 14096 13719 14148 13728
rect 14096 13685 14105 13719
rect 14105 13685 14139 13719
rect 14139 13685 14148 13719
rect 14096 13676 14148 13685
rect 14832 13676 14884 13728
rect 15200 13719 15252 13728
rect 15200 13685 15209 13719
rect 15209 13685 15243 13719
rect 15243 13685 15252 13719
rect 15200 13676 15252 13685
rect 15936 13676 15988 13728
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 19022 13574 19074 13626
rect 19086 13574 19138 13626
rect 19150 13574 19202 13626
rect 19214 13574 19266 13626
rect 19278 13574 19330 13626
rect 4068 13472 4120 13524
rect 5632 13515 5684 13524
rect 5632 13481 5641 13515
rect 5641 13481 5675 13515
rect 5675 13481 5684 13515
rect 5632 13472 5684 13481
rect 8576 13472 8628 13524
rect 5356 13404 5408 13456
rect 4160 13268 4212 13320
rect 6828 13336 6880 13388
rect 7932 13379 7984 13388
rect 7932 13345 7941 13379
rect 7941 13345 7975 13379
rect 7975 13345 7984 13379
rect 7932 13336 7984 13345
rect 8208 13379 8260 13388
rect 8208 13345 8217 13379
rect 8217 13345 8251 13379
rect 8251 13345 8260 13379
rect 8208 13336 8260 13345
rect 8392 13379 8444 13388
rect 8392 13345 8401 13379
rect 8401 13345 8435 13379
rect 8435 13345 8444 13379
rect 8392 13336 8444 13345
rect 17040 13472 17092 13524
rect 7380 13268 7432 13320
rect 8300 13268 8352 13320
rect 9772 13336 9824 13388
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 10048 13311 10100 13320
rect 10048 13277 10057 13311
rect 10057 13277 10091 13311
rect 10091 13277 10100 13311
rect 10048 13268 10100 13277
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 10968 13336 11020 13388
rect 16212 13404 16264 13456
rect 19800 13404 19852 13456
rect 11428 13336 11480 13388
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 14556 13379 14608 13388
rect 14556 13345 14565 13379
rect 14565 13345 14599 13379
rect 14599 13345 14608 13379
rect 14556 13336 14608 13345
rect 15108 13336 15160 13388
rect 16120 13379 16172 13388
rect 16120 13345 16129 13379
rect 16129 13345 16163 13379
rect 16163 13345 16172 13379
rect 16120 13336 16172 13345
rect 11060 13311 11112 13320
rect 11060 13277 11069 13311
rect 11069 13277 11103 13311
rect 11103 13277 11112 13311
rect 11060 13268 11112 13277
rect 11796 13268 11848 13320
rect 19340 13379 19392 13388
rect 19340 13345 19349 13379
rect 19349 13345 19383 13379
rect 19383 13345 19392 13379
rect 19340 13336 19392 13345
rect 20536 13472 20588 13524
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 20444 13336 20496 13388
rect 21180 13404 21232 13456
rect 21272 13336 21324 13388
rect 12900 13200 12952 13252
rect 18788 13200 18840 13252
rect 4528 13132 4580 13184
rect 8300 13175 8352 13184
rect 8300 13141 8309 13175
rect 8309 13141 8343 13175
rect 8343 13141 8352 13175
rect 8300 13132 8352 13141
rect 9864 13175 9916 13184
rect 9864 13141 9873 13175
rect 9873 13141 9907 13175
rect 9907 13141 9916 13175
rect 9864 13132 9916 13141
rect 11520 13175 11572 13184
rect 11520 13141 11529 13175
rect 11529 13141 11563 13175
rect 11563 13141 11572 13175
rect 11520 13132 11572 13141
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 17592 13132 17644 13184
rect 18420 13132 18472 13184
rect 20812 13200 20864 13252
rect 20076 13175 20128 13184
rect 20076 13141 20085 13175
rect 20085 13141 20119 13175
rect 20119 13141 20128 13175
rect 20076 13132 20128 13141
rect 21272 13175 21324 13184
rect 21272 13141 21281 13175
rect 21281 13141 21315 13175
rect 21315 13141 21324 13175
rect 21272 13132 21324 13141
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 8300 12928 8352 12980
rect 10324 12928 10376 12980
rect 15108 12928 15160 12980
rect 16028 12928 16080 12980
rect 17684 12928 17736 12980
rect 20720 12928 20772 12980
rect 21456 12928 21508 12980
rect 4252 12767 4304 12776
rect 4252 12733 4261 12767
rect 4261 12733 4295 12767
rect 4295 12733 4304 12767
rect 4252 12724 4304 12733
rect 4528 12767 4580 12776
rect 4528 12733 4537 12767
rect 4537 12733 4571 12767
rect 4571 12733 4580 12767
rect 4528 12724 4580 12733
rect 15292 12860 15344 12912
rect 7472 12656 7524 12708
rect 9404 12656 9456 12708
rect 9956 12656 10008 12708
rect 10784 12767 10836 12776
rect 10784 12733 10793 12767
rect 10793 12733 10827 12767
rect 10827 12733 10836 12767
rect 10784 12724 10836 12733
rect 14096 12792 14148 12844
rect 11336 12656 11388 12708
rect 13912 12724 13964 12776
rect 15476 12792 15528 12844
rect 15844 12835 15896 12844
rect 15844 12801 15853 12835
rect 15853 12801 15887 12835
rect 15887 12801 15896 12835
rect 15844 12792 15896 12801
rect 15108 12724 15160 12776
rect 15200 12724 15252 12776
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 19432 12792 19484 12844
rect 16948 12724 17000 12776
rect 17592 12767 17644 12776
rect 17592 12733 17601 12767
rect 17601 12733 17635 12767
rect 17635 12733 17644 12767
rect 17592 12724 17644 12733
rect 17776 12724 17828 12776
rect 19340 12724 19392 12776
rect 20996 12903 21048 12912
rect 20996 12869 21005 12903
rect 21005 12869 21039 12903
rect 21039 12869 21048 12903
rect 20996 12860 21048 12869
rect 22100 12860 22152 12912
rect 22468 12792 22520 12844
rect 22652 12835 22704 12844
rect 22652 12801 22661 12835
rect 22661 12801 22695 12835
rect 22695 12801 22704 12835
rect 22652 12792 22704 12801
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 21180 12724 21232 12776
rect 21456 12767 21508 12776
rect 21456 12733 21465 12767
rect 21465 12733 21499 12767
rect 21499 12733 21508 12767
rect 21456 12724 21508 12733
rect 21732 12724 21784 12776
rect 22744 12767 22796 12776
rect 22744 12733 22753 12767
rect 22753 12733 22787 12767
rect 22787 12733 22796 12767
rect 22744 12724 22796 12733
rect 5908 12631 5960 12640
rect 5908 12597 5917 12631
rect 5917 12597 5951 12631
rect 5951 12597 5960 12631
rect 5908 12588 5960 12597
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 8484 12588 8536 12640
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 14372 12631 14424 12640
rect 14372 12597 14381 12631
rect 14381 12597 14415 12631
rect 14415 12597 14424 12631
rect 14372 12588 14424 12597
rect 14832 12699 14884 12708
rect 14832 12665 14841 12699
rect 14841 12665 14875 12699
rect 14875 12665 14884 12699
rect 14832 12656 14884 12665
rect 17224 12656 17276 12708
rect 21364 12656 21416 12708
rect 20720 12588 20772 12640
rect 21088 12631 21140 12640
rect 21088 12597 21097 12631
rect 21097 12597 21131 12631
rect 21131 12597 21140 12631
rect 21088 12588 21140 12597
rect 22192 12588 22244 12640
rect 19022 12486 19074 12538
rect 19086 12486 19138 12538
rect 19150 12486 19202 12538
rect 19214 12486 19266 12538
rect 19278 12486 19330 12538
rect 4252 12384 4304 12436
rect 5264 12427 5316 12436
rect 5264 12393 5273 12427
rect 5273 12393 5307 12427
rect 5307 12393 5316 12427
rect 5264 12384 5316 12393
rect 5908 12384 5960 12436
rect 7472 12427 7524 12436
rect 7472 12393 7481 12427
rect 7481 12393 7515 12427
rect 7515 12393 7524 12427
rect 7472 12384 7524 12393
rect 7840 12384 7892 12436
rect 8392 12384 8444 12436
rect 10784 12427 10836 12436
rect 10784 12393 10793 12427
rect 10793 12393 10827 12427
rect 10827 12393 10836 12427
rect 10784 12384 10836 12393
rect 12900 12427 12952 12436
rect 12900 12393 12909 12427
rect 12909 12393 12943 12427
rect 12943 12393 12952 12427
rect 12900 12384 12952 12393
rect 5540 12316 5592 12368
rect 8484 12316 8536 12368
rect 9864 12316 9916 12368
rect 9956 12316 10008 12368
rect 11520 12316 11572 12368
rect 12348 12316 12400 12368
rect 13728 12384 13780 12436
rect 14372 12384 14424 12436
rect 20352 12384 20404 12436
rect 16304 12316 16356 12368
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 7932 12291 7984 12300
rect 7932 12257 7941 12291
rect 7941 12257 7975 12291
rect 7975 12257 7984 12291
rect 7932 12248 7984 12257
rect 13452 12291 13504 12300
rect 13452 12257 13461 12291
rect 13461 12257 13495 12291
rect 13495 12257 13504 12291
rect 13452 12248 13504 12257
rect 13820 12248 13872 12300
rect 15384 12291 15436 12300
rect 15384 12257 15393 12291
rect 15393 12257 15427 12291
rect 15427 12257 15436 12291
rect 15384 12248 15436 12257
rect 16948 12291 17000 12300
rect 16948 12257 16957 12291
rect 16957 12257 16991 12291
rect 16991 12257 17000 12291
rect 16948 12248 17000 12257
rect 17224 12291 17276 12300
rect 17224 12257 17233 12291
rect 17233 12257 17267 12291
rect 17267 12257 17276 12291
rect 17224 12248 17276 12257
rect 17776 12248 17828 12300
rect 21088 12316 21140 12368
rect 21916 12384 21968 12436
rect 18788 12248 18840 12300
rect 20812 12291 20864 12300
rect 20812 12257 20821 12291
rect 20821 12257 20855 12291
rect 20855 12257 20864 12291
rect 20812 12248 20864 12257
rect 20904 12248 20956 12300
rect 8208 12112 8260 12164
rect 9588 12044 9640 12096
rect 10968 12087 11020 12096
rect 10968 12053 10977 12087
rect 10977 12053 11011 12087
rect 11011 12053 11020 12087
rect 10968 12044 11020 12053
rect 12440 12087 12492 12096
rect 12440 12053 12449 12087
rect 12449 12053 12483 12087
rect 12483 12053 12492 12087
rect 12440 12044 12492 12053
rect 13636 12044 13688 12096
rect 16856 12180 16908 12232
rect 17684 12180 17736 12232
rect 20996 12180 21048 12232
rect 22192 12248 22244 12300
rect 22284 12291 22336 12300
rect 22284 12257 22293 12291
rect 22293 12257 22327 12291
rect 22327 12257 22336 12291
rect 22284 12248 22336 12257
rect 23296 12248 23348 12300
rect 14372 12044 14424 12096
rect 15108 12087 15160 12096
rect 15108 12053 15117 12087
rect 15117 12053 15151 12087
rect 15151 12053 15160 12087
rect 15108 12044 15160 12053
rect 15200 12087 15252 12096
rect 15200 12053 15209 12087
rect 15209 12053 15243 12087
rect 15243 12053 15252 12087
rect 15200 12044 15252 12053
rect 18236 12087 18288 12096
rect 18236 12053 18245 12087
rect 18245 12053 18279 12087
rect 18279 12053 18288 12087
rect 18236 12044 18288 12053
rect 21272 12087 21324 12096
rect 21272 12053 21281 12087
rect 21281 12053 21315 12087
rect 21315 12053 21324 12087
rect 21272 12044 21324 12053
rect 22100 12087 22152 12096
rect 22100 12053 22109 12087
rect 22109 12053 22143 12087
rect 22143 12053 22152 12087
rect 22100 12044 22152 12053
rect 22376 12087 22428 12096
rect 22376 12053 22385 12087
rect 22385 12053 22419 12087
rect 22419 12053 22428 12087
rect 22376 12044 22428 12053
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 5724 11883 5776 11892
rect 5724 11849 5733 11883
rect 5733 11849 5767 11883
rect 5767 11849 5776 11883
rect 5724 11840 5776 11849
rect 11060 11840 11112 11892
rect 12440 11840 12492 11892
rect 13912 11840 13964 11892
rect 15108 11883 15160 11892
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 15200 11840 15252 11892
rect 18236 11840 18288 11892
rect 20904 11840 20956 11892
rect 21456 11840 21508 11892
rect 5540 11772 5592 11824
rect 10968 11704 11020 11756
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 6000 11679 6052 11688
rect 6000 11645 6009 11679
rect 6009 11645 6043 11679
rect 6043 11645 6052 11679
rect 6000 11636 6052 11645
rect 6460 11636 6512 11688
rect 7656 11636 7708 11688
rect 11336 11679 11388 11688
rect 11336 11645 11345 11679
rect 11345 11645 11379 11679
rect 11379 11645 11388 11679
rect 11336 11636 11388 11645
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 15936 11704 15988 11756
rect 17224 11772 17276 11824
rect 16304 11704 16356 11756
rect 16396 11747 16448 11756
rect 16396 11713 16405 11747
rect 16405 11713 16439 11747
rect 16439 11713 16448 11747
rect 16396 11704 16448 11713
rect 8576 11568 8628 11620
rect 13820 11568 13872 11620
rect 15016 11568 15068 11620
rect 5816 11500 5868 11552
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 7196 11500 7248 11552
rect 8668 11500 8720 11552
rect 11980 11543 12032 11552
rect 11980 11509 11989 11543
rect 11989 11509 12023 11543
rect 12023 11509 12032 11543
rect 11980 11500 12032 11509
rect 14556 11500 14608 11552
rect 14740 11500 14792 11552
rect 16856 11636 16908 11688
rect 16948 11636 17000 11688
rect 19432 11747 19484 11756
rect 19432 11713 19441 11747
rect 19441 11713 19475 11747
rect 19475 11713 19484 11747
rect 19432 11704 19484 11713
rect 18788 11568 18840 11620
rect 19524 11679 19576 11688
rect 19524 11645 19533 11679
rect 19533 11645 19567 11679
rect 19567 11645 19576 11679
rect 19524 11636 19576 11645
rect 20260 11679 20312 11688
rect 20260 11645 20269 11679
rect 20269 11645 20303 11679
rect 20303 11645 20312 11679
rect 20260 11636 20312 11645
rect 22560 11636 22612 11688
rect 19984 11611 20036 11620
rect 19984 11577 19993 11611
rect 19993 11577 20027 11611
rect 20027 11577 20036 11611
rect 19984 11568 20036 11577
rect 22284 11568 22336 11620
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 20996 11500 21048 11552
rect 22376 11500 22428 11552
rect 19022 11398 19074 11450
rect 19086 11398 19138 11450
rect 19150 11398 19202 11450
rect 19214 11398 19266 11450
rect 19278 11398 19330 11450
rect 6184 11296 6236 11348
rect 5448 11228 5500 11280
rect 7288 11339 7340 11348
rect 7288 11305 7313 11339
rect 7313 11305 7340 11339
rect 7288 11296 7340 11305
rect 9680 11296 9732 11348
rect 5724 11160 5776 11212
rect 7564 11228 7616 11280
rect 5816 11092 5868 11144
rect 5724 11024 5776 11076
rect 5540 10999 5592 11008
rect 5540 10965 5549 10999
rect 5549 10965 5583 10999
rect 5583 10965 5592 10999
rect 5540 10956 5592 10965
rect 5908 10956 5960 11008
rect 6092 11024 6144 11076
rect 7656 11203 7708 11212
rect 7656 11169 7665 11203
rect 7665 11169 7699 11203
rect 7699 11169 7708 11203
rect 7656 11160 7708 11169
rect 8208 11160 8260 11212
rect 6276 10956 6328 11008
rect 6552 10999 6604 11008
rect 6552 10965 6561 10999
rect 6561 10965 6595 10999
rect 6595 10965 6604 10999
rect 6552 10956 6604 10965
rect 7196 10956 7248 11008
rect 8576 11271 8628 11280
rect 8576 11237 8585 11271
rect 8585 11237 8619 11271
rect 8619 11237 8628 11271
rect 8576 11228 8628 11237
rect 8484 11203 8536 11212
rect 8484 11169 8493 11203
rect 8493 11169 8527 11203
rect 8527 11169 8536 11203
rect 8484 11160 8536 11169
rect 10784 11160 10836 11212
rect 11980 11296 12032 11348
rect 12348 11296 12400 11348
rect 16304 11296 16356 11348
rect 16948 11296 17000 11348
rect 19984 11296 20036 11348
rect 20996 11296 21048 11348
rect 22100 11296 22152 11348
rect 9864 11024 9916 11076
rect 10968 11024 11020 11076
rect 7840 10956 7892 11008
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 8484 10956 8536 11008
rect 8668 10956 8720 11008
rect 10048 10956 10100 11008
rect 12624 11160 12676 11212
rect 13912 11160 13964 11212
rect 14096 11160 14148 11212
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 14280 11160 14332 11212
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 15292 11160 15344 11212
rect 16396 11160 16448 11212
rect 18880 11203 18932 11212
rect 18880 11169 18889 11203
rect 18889 11169 18923 11203
rect 18923 11169 18932 11203
rect 18880 11160 18932 11169
rect 15016 11135 15068 11144
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15016 11092 15068 11101
rect 19892 11160 19944 11212
rect 21364 11228 21416 11280
rect 22008 11228 22060 11280
rect 20904 11092 20956 11144
rect 15108 11024 15160 11076
rect 20536 11067 20588 11076
rect 20536 11033 20545 11067
rect 20545 11033 20579 11067
rect 20579 11033 20588 11067
rect 20536 11024 20588 11033
rect 11888 10956 11940 11008
rect 12256 10956 12308 11008
rect 14004 10956 14056 11008
rect 14188 10999 14240 11008
rect 14188 10965 14197 10999
rect 14197 10965 14231 10999
rect 14231 10965 14240 10999
rect 14188 10956 14240 10965
rect 16212 10999 16264 11008
rect 16212 10965 16221 10999
rect 16221 10965 16255 10999
rect 16255 10965 16264 10999
rect 16212 10956 16264 10965
rect 16764 10999 16816 11008
rect 16764 10965 16773 10999
rect 16773 10965 16807 10999
rect 16807 10965 16816 10999
rect 16764 10956 16816 10965
rect 19616 10956 19668 11008
rect 20996 10956 21048 11008
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 5448 10752 5500 10804
rect 6184 10752 6236 10804
rect 6276 10795 6328 10804
rect 6276 10761 6285 10795
rect 6285 10761 6319 10795
rect 6319 10761 6328 10795
rect 6276 10752 6328 10761
rect 9680 10752 9732 10804
rect 10968 10752 11020 10804
rect 20260 10752 20312 10804
rect 20536 10752 20588 10804
rect 20904 10795 20956 10804
rect 20904 10761 20913 10795
rect 20913 10761 20947 10795
rect 20947 10761 20956 10795
rect 20904 10752 20956 10761
rect 20996 10752 21048 10804
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 6644 10591 6696 10600
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 7288 10548 7340 10600
rect 7840 10684 7892 10736
rect 8392 10684 8444 10736
rect 8208 10616 8260 10668
rect 8668 10659 8720 10668
rect 8668 10625 8677 10659
rect 8677 10625 8711 10659
rect 8711 10625 8720 10659
rect 8668 10616 8720 10625
rect 5540 10412 5592 10464
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 5632 10412 5684 10421
rect 7196 10412 7248 10464
rect 7748 10523 7800 10532
rect 7748 10489 7757 10523
rect 7757 10489 7791 10523
rect 7791 10489 7800 10523
rect 7748 10480 7800 10489
rect 10600 10684 10652 10736
rect 9036 10523 9088 10532
rect 9036 10489 9045 10523
rect 9045 10489 9079 10523
rect 9079 10489 9088 10523
rect 9036 10480 9088 10489
rect 9864 10591 9916 10600
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 10048 10591 10100 10600
rect 10048 10557 10057 10591
rect 10057 10557 10091 10591
rect 10091 10557 10100 10591
rect 10048 10548 10100 10557
rect 10692 10659 10744 10668
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 9680 10480 9732 10532
rect 10600 10548 10652 10600
rect 10968 10548 11020 10600
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 12624 10591 12676 10600
rect 12624 10557 12633 10591
rect 12633 10557 12667 10591
rect 12667 10557 12676 10591
rect 12624 10548 12676 10557
rect 14188 10616 14240 10668
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 14280 10591 14332 10600
rect 14280 10557 14289 10591
rect 14289 10557 14323 10591
rect 14323 10557 14332 10591
rect 14280 10548 14332 10557
rect 16212 10616 16264 10668
rect 16764 10659 16816 10668
rect 16764 10625 16773 10659
rect 16773 10625 16807 10659
rect 16807 10625 16816 10659
rect 16764 10616 16816 10625
rect 16856 10616 16908 10668
rect 20720 10684 20772 10736
rect 21548 10684 21600 10736
rect 22284 10795 22336 10804
rect 22284 10761 22293 10795
rect 22293 10761 22327 10795
rect 22327 10761 22336 10795
rect 22284 10752 22336 10761
rect 14096 10480 14148 10532
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 16672 10591 16724 10600
rect 16672 10557 16681 10591
rect 16681 10557 16715 10591
rect 16715 10557 16724 10591
rect 16672 10548 16724 10557
rect 17316 10591 17368 10600
rect 17316 10557 17325 10591
rect 17325 10557 17359 10591
rect 17359 10557 17368 10591
rect 17316 10548 17368 10557
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 9404 10412 9456 10464
rect 9496 10455 9548 10464
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 9772 10455 9824 10464
rect 9772 10421 9781 10455
rect 9781 10421 9815 10455
rect 9815 10421 9824 10455
rect 9772 10412 9824 10421
rect 11060 10412 11112 10464
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 13912 10412 13964 10464
rect 14832 10455 14884 10464
rect 14832 10421 14841 10455
rect 14841 10421 14875 10455
rect 14875 10421 14884 10455
rect 14832 10412 14884 10421
rect 20904 10523 20956 10532
rect 20904 10489 20913 10523
rect 20913 10489 20947 10523
rect 20947 10489 20956 10523
rect 20904 10480 20956 10489
rect 21456 10548 21508 10600
rect 22100 10591 22152 10600
rect 22100 10557 22109 10591
rect 22109 10557 22143 10591
rect 22143 10557 22152 10591
rect 22100 10548 22152 10557
rect 22008 10523 22060 10532
rect 22008 10489 22017 10523
rect 22017 10489 22051 10523
rect 22051 10489 22060 10523
rect 22008 10480 22060 10489
rect 20628 10412 20680 10464
rect 21364 10412 21416 10464
rect 19022 10310 19074 10362
rect 19086 10310 19138 10362
rect 19150 10310 19202 10362
rect 19214 10310 19266 10362
rect 19278 10310 19330 10362
rect 6644 10208 6696 10260
rect 5264 10183 5316 10192
rect 5264 10149 5273 10183
rect 5273 10149 5307 10183
rect 5307 10149 5316 10183
rect 5264 10140 5316 10149
rect 5632 10072 5684 10124
rect 6092 10004 6144 10056
rect 8392 10208 8444 10260
rect 9036 10208 9088 10260
rect 9404 10251 9456 10260
rect 9404 10217 9413 10251
rect 9413 10217 9447 10251
rect 9447 10217 9456 10251
rect 9404 10208 9456 10217
rect 9680 10208 9732 10260
rect 9772 10208 9824 10260
rect 10692 10208 10744 10260
rect 11244 10208 11296 10260
rect 18052 10208 18104 10260
rect 20904 10208 20956 10260
rect 8392 10115 8444 10124
rect 8392 10081 8401 10115
rect 8401 10081 8435 10115
rect 8435 10081 8444 10115
rect 8392 10072 8444 10081
rect 8576 10072 8628 10124
rect 10508 10072 10560 10124
rect 22744 10140 22796 10192
rect 14096 10072 14148 10124
rect 14464 10115 14516 10124
rect 14464 10081 14473 10115
rect 14473 10081 14507 10115
rect 14507 10081 14516 10115
rect 14464 10072 14516 10081
rect 19616 10115 19668 10124
rect 19616 10081 19625 10115
rect 19625 10081 19659 10115
rect 19659 10081 19668 10115
rect 19616 10072 19668 10081
rect 19708 10115 19760 10124
rect 19708 10081 19717 10115
rect 19717 10081 19751 10115
rect 19751 10081 19760 10115
rect 19708 10072 19760 10081
rect 19892 10115 19944 10124
rect 19892 10081 19901 10115
rect 19901 10081 19935 10115
rect 19935 10081 19944 10115
rect 19892 10072 19944 10081
rect 21364 10072 21416 10124
rect 21548 10115 21600 10124
rect 21548 10081 21557 10115
rect 21557 10081 21591 10115
rect 21591 10081 21600 10115
rect 21548 10072 21600 10081
rect 21732 10115 21784 10124
rect 21732 10081 21741 10115
rect 21741 10081 21775 10115
rect 21775 10081 21784 10115
rect 21732 10072 21784 10081
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 5632 9979 5684 9988
rect 5632 9945 5641 9979
rect 5641 9945 5675 9979
rect 5675 9945 5684 9979
rect 5632 9936 5684 9945
rect 6276 9936 6328 9988
rect 9496 9936 9548 9988
rect 11704 9936 11756 9988
rect 4252 9868 4304 9920
rect 6552 9868 6604 9920
rect 10600 9911 10652 9920
rect 10600 9877 10609 9911
rect 10609 9877 10643 9911
rect 10643 9877 10652 9911
rect 10600 9868 10652 9877
rect 11152 9911 11204 9920
rect 11152 9877 11161 9911
rect 11161 9877 11195 9911
rect 11195 9877 11204 9911
rect 11152 9868 11204 9877
rect 14188 9911 14240 9920
rect 14188 9877 14197 9911
rect 14197 9877 14231 9911
rect 14231 9877 14240 9911
rect 14188 9868 14240 9877
rect 18880 9868 18932 9920
rect 19248 9868 19300 9920
rect 20904 10004 20956 10056
rect 20536 9936 20588 9988
rect 20628 9868 20680 9920
rect 21364 9911 21416 9920
rect 21364 9877 21373 9911
rect 21373 9877 21407 9911
rect 21407 9877 21416 9911
rect 21364 9868 21416 9877
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 5724 9707 5776 9716
rect 5724 9673 5733 9707
rect 5733 9673 5767 9707
rect 5767 9673 5776 9707
rect 5724 9664 5776 9673
rect 6552 9707 6604 9716
rect 6552 9673 6561 9707
rect 6561 9673 6595 9707
rect 6595 9673 6604 9707
rect 6552 9664 6604 9673
rect 5632 9596 5684 9648
rect 10600 9664 10652 9716
rect 14188 9664 14240 9716
rect 14280 9707 14332 9716
rect 14280 9673 14289 9707
rect 14289 9673 14323 9707
rect 14323 9673 14332 9707
rect 14280 9664 14332 9673
rect 14464 9664 14516 9716
rect 4252 9460 4304 9512
rect 4344 9503 4396 9512
rect 4344 9469 4353 9503
rect 4353 9469 4387 9503
rect 4387 9469 4396 9503
rect 4344 9460 4396 9469
rect 5724 9460 5776 9512
rect 6184 9460 6236 9512
rect 11060 9528 11112 9580
rect 11152 9528 11204 9580
rect 18236 9596 18288 9648
rect 12808 9528 12860 9580
rect 14832 9528 14884 9580
rect 19708 9664 19760 9716
rect 19892 9664 19944 9716
rect 20720 9664 20772 9716
rect 20812 9664 20864 9716
rect 21732 9664 21784 9716
rect 20076 9639 20128 9648
rect 20076 9605 20085 9639
rect 20085 9605 20119 9639
rect 20119 9605 20128 9639
rect 20076 9596 20128 9605
rect 7012 9503 7064 9512
rect 7012 9469 7021 9503
rect 7021 9469 7055 9503
rect 7055 9469 7064 9503
rect 7012 9460 7064 9469
rect 10968 9503 11020 9512
rect 10968 9469 10977 9503
rect 10977 9469 11011 9503
rect 11011 9469 11020 9503
rect 10968 9460 11020 9469
rect 6276 9392 6328 9444
rect 11060 9392 11112 9444
rect 11704 9460 11756 9512
rect 13728 9503 13780 9512
rect 13728 9469 13737 9503
rect 13737 9469 13771 9503
rect 13771 9469 13780 9503
rect 13728 9460 13780 9469
rect 14188 9460 14240 9512
rect 16856 9460 16908 9512
rect 5540 9324 5592 9376
rect 5724 9324 5776 9376
rect 6092 9324 6144 9376
rect 6460 9324 6512 9376
rect 7012 9324 7064 9376
rect 17684 9392 17736 9444
rect 18696 9460 18748 9512
rect 18788 9503 18840 9512
rect 18788 9469 18797 9503
rect 18797 9469 18831 9503
rect 18831 9469 18840 9503
rect 18788 9460 18840 9469
rect 16488 9367 16540 9376
rect 16488 9333 16497 9367
rect 16497 9333 16531 9367
rect 16531 9333 16540 9367
rect 16488 9324 16540 9333
rect 18144 9435 18196 9444
rect 18144 9401 18153 9435
rect 18153 9401 18187 9435
rect 18187 9401 18196 9435
rect 19248 9528 19300 9580
rect 19340 9460 19392 9512
rect 18144 9392 18196 9401
rect 19524 9460 19576 9512
rect 22560 9596 22612 9648
rect 20168 9460 20220 9512
rect 20352 9392 20404 9444
rect 19708 9324 19760 9376
rect 20168 9324 20220 9376
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 21088 9460 21140 9512
rect 21364 9392 21416 9444
rect 20720 9324 20772 9376
rect 20812 9324 20864 9376
rect 20904 9367 20956 9376
rect 20904 9333 20913 9367
rect 20913 9333 20947 9367
rect 20947 9333 20956 9367
rect 20904 9324 20956 9333
rect 22100 9324 22152 9376
rect 19022 9222 19074 9274
rect 19086 9222 19138 9274
rect 19150 9222 19202 9274
rect 19214 9222 19266 9274
rect 19278 9222 19330 9274
rect 4344 9120 4396 9172
rect 6184 9120 6236 9172
rect 6460 9120 6512 9172
rect 8760 9120 8812 9172
rect 14096 9120 14148 9172
rect 16488 9120 16540 9172
rect 17316 9120 17368 9172
rect 17960 9120 18012 9172
rect 18236 9120 18288 9172
rect 18696 9120 18748 9172
rect 7104 9052 7156 9104
rect 4896 8984 4948 9036
rect 6368 8984 6420 9036
rect 7748 9052 7800 9104
rect 14924 9052 14976 9104
rect 18788 9052 18840 9104
rect 19708 9052 19760 9104
rect 19800 9095 19852 9104
rect 19800 9061 19809 9095
rect 19809 9061 19843 9095
rect 19843 9061 19852 9095
rect 19800 9052 19852 9061
rect 16856 8984 16908 9036
rect 20076 8984 20128 9036
rect 13912 8959 13964 8968
rect 13912 8925 13921 8959
rect 13921 8925 13955 8959
rect 13955 8925 13964 8959
rect 13912 8916 13964 8925
rect 5172 8780 5224 8832
rect 5540 8780 5592 8832
rect 5816 8780 5868 8832
rect 7564 8780 7616 8832
rect 7932 8780 7984 8832
rect 14556 8848 14608 8900
rect 18144 8959 18196 8968
rect 18144 8925 18153 8959
rect 18153 8925 18187 8959
rect 18187 8925 18196 8959
rect 18144 8916 18196 8925
rect 19432 8916 19484 8968
rect 19524 8916 19576 8968
rect 19708 8916 19760 8968
rect 20352 9027 20404 9036
rect 20352 8993 20361 9027
rect 20361 8993 20395 9027
rect 20395 8993 20404 9027
rect 20352 8984 20404 8993
rect 20904 9120 20956 9172
rect 21088 9120 21140 9172
rect 21272 9120 21324 9172
rect 22560 9120 22612 9172
rect 22744 9120 22796 9172
rect 22008 8984 22060 9036
rect 8116 8780 8168 8832
rect 8576 8780 8628 8832
rect 9588 8780 9640 8832
rect 14464 8780 14516 8832
rect 16120 8780 16172 8832
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 19984 8848 20036 8900
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 20168 8780 20220 8832
rect 20628 8780 20680 8832
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 5080 8576 5132 8628
rect 5356 8619 5408 8628
rect 5356 8585 5365 8619
rect 5365 8585 5399 8619
rect 5399 8585 5408 8619
rect 5356 8576 5408 8585
rect 5632 8576 5684 8628
rect 6184 8576 6236 8628
rect 6368 8576 6420 8628
rect 5724 8508 5776 8560
rect 5816 8508 5868 8560
rect 5080 8372 5132 8424
rect 7288 8551 7340 8560
rect 7288 8517 7297 8551
rect 7297 8517 7331 8551
rect 7331 8517 7340 8551
rect 7288 8508 7340 8517
rect 7564 8508 7616 8560
rect 7932 8576 7984 8628
rect 10140 8576 10192 8628
rect 8300 8508 8352 8560
rect 5172 8236 5224 8288
rect 6460 8415 6512 8424
rect 6460 8381 6469 8415
rect 6469 8381 6503 8415
rect 6503 8381 6512 8415
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 8392 8440 8444 8492
rect 6460 8372 6512 8381
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 8760 8440 8812 8492
rect 10140 8440 10192 8492
rect 9036 8372 9088 8424
rect 10784 8440 10836 8492
rect 12532 8508 12584 8560
rect 13728 8508 13780 8560
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 10968 8372 11020 8424
rect 13636 8440 13688 8492
rect 7748 8236 7800 8288
rect 10692 8304 10744 8356
rect 11244 8372 11296 8424
rect 13176 8372 13228 8424
rect 14740 8576 14792 8628
rect 16672 8576 16724 8628
rect 17224 8619 17276 8628
rect 17224 8585 17233 8619
rect 17233 8585 17267 8619
rect 17267 8585 17276 8619
rect 17224 8576 17276 8585
rect 17684 8619 17736 8628
rect 17684 8585 17693 8619
rect 17693 8585 17727 8619
rect 17727 8585 17736 8619
rect 17684 8576 17736 8585
rect 18052 8576 18104 8628
rect 18144 8576 18196 8628
rect 18696 8576 18748 8628
rect 19616 8576 19668 8628
rect 19708 8576 19760 8628
rect 20628 8619 20680 8628
rect 20628 8585 20637 8619
rect 20637 8585 20671 8619
rect 20671 8585 20680 8619
rect 20628 8576 20680 8585
rect 21824 8576 21876 8628
rect 14004 8508 14056 8560
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 15660 8551 15712 8560
rect 15660 8517 15669 8551
rect 15669 8517 15703 8551
rect 15703 8517 15712 8551
rect 15660 8508 15712 8517
rect 16028 8508 16080 8560
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 14832 8415 14884 8424
rect 14832 8381 14841 8415
rect 14841 8381 14875 8415
rect 14875 8381 14884 8415
rect 14832 8372 14884 8381
rect 10232 8279 10284 8288
rect 10232 8245 10241 8279
rect 10241 8245 10275 8279
rect 10275 8245 10284 8279
rect 10232 8236 10284 8245
rect 10508 8236 10560 8288
rect 11060 8236 11112 8288
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 11612 8236 11664 8288
rect 12716 8279 12768 8288
rect 12716 8245 12725 8279
rect 12725 8245 12759 8279
rect 12759 8245 12768 8279
rect 12716 8236 12768 8245
rect 13728 8279 13780 8288
rect 13728 8245 13737 8279
rect 13737 8245 13771 8279
rect 13771 8245 13780 8279
rect 13728 8236 13780 8245
rect 14372 8279 14424 8288
rect 14372 8245 14381 8279
rect 14381 8245 14415 8279
rect 14415 8245 14424 8279
rect 14372 8236 14424 8245
rect 14648 8347 14700 8356
rect 14648 8313 14657 8347
rect 14657 8313 14691 8347
rect 14691 8313 14700 8347
rect 14648 8304 14700 8313
rect 15108 8415 15160 8424
rect 15108 8381 15117 8415
rect 15117 8381 15151 8415
rect 15151 8381 15160 8415
rect 15108 8372 15160 8381
rect 16672 8440 16724 8492
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 17316 8440 17368 8492
rect 17868 8508 17920 8560
rect 18696 8415 18748 8424
rect 18696 8381 18705 8415
rect 18705 8381 18739 8415
rect 18739 8381 18748 8415
rect 18696 8372 18748 8381
rect 20812 8508 20864 8560
rect 20536 8372 20588 8424
rect 21548 8483 21600 8492
rect 21548 8449 21557 8483
rect 21557 8449 21591 8483
rect 21591 8449 21600 8483
rect 21548 8440 21600 8449
rect 21732 8483 21784 8492
rect 21732 8449 21741 8483
rect 21741 8449 21775 8483
rect 21775 8449 21784 8483
rect 21732 8440 21784 8449
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 14924 8236 14976 8288
rect 15292 8236 15344 8288
rect 16028 8304 16080 8356
rect 17408 8347 17460 8356
rect 17408 8313 17417 8347
rect 17417 8313 17451 8347
rect 17451 8313 17460 8347
rect 17408 8304 17460 8313
rect 22100 8304 22152 8356
rect 22744 8304 22796 8356
rect 17684 8236 17736 8288
rect 21088 8279 21140 8288
rect 21088 8245 21097 8279
rect 21097 8245 21131 8279
rect 21131 8245 21140 8279
rect 21088 8236 21140 8245
rect 22008 8279 22060 8288
rect 22008 8245 22017 8279
rect 22017 8245 22051 8279
rect 22051 8245 22060 8279
rect 22008 8236 22060 8245
rect 22652 8279 22704 8288
rect 22652 8245 22661 8279
rect 22661 8245 22695 8279
rect 22695 8245 22704 8279
rect 22652 8236 22704 8245
rect 19022 8134 19074 8186
rect 19086 8134 19138 8186
rect 19150 8134 19202 8186
rect 19214 8134 19266 8186
rect 19278 8134 19330 8186
rect 7748 8075 7800 8084
rect 7748 8041 7757 8075
rect 7757 8041 7791 8075
rect 7791 8041 7800 8075
rect 7748 8032 7800 8041
rect 8392 8032 8444 8084
rect 10968 8075 11020 8084
rect 10968 8041 10977 8075
rect 10977 8041 11011 8075
rect 11011 8041 11020 8075
rect 10968 8032 11020 8041
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 12716 8032 12768 8084
rect 13176 8032 13228 8084
rect 13268 8032 13320 8084
rect 13728 8032 13780 8084
rect 14188 8075 14240 8084
rect 14188 8041 14197 8075
rect 14197 8041 14231 8075
rect 14231 8041 14240 8075
rect 14188 8032 14240 8041
rect 7288 7964 7340 8016
rect 5908 7896 5960 7948
rect 7104 7896 7156 7948
rect 8944 7939 8996 7948
rect 9588 7964 9640 8016
rect 10692 8007 10744 8016
rect 10692 7973 10701 8007
rect 10701 7973 10735 8007
rect 10735 7973 10744 8007
rect 10692 7964 10744 7973
rect 10784 7964 10836 8016
rect 8944 7905 8962 7939
rect 8962 7905 8996 7939
rect 8944 7896 8996 7905
rect 9864 7803 9916 7812
rect 9864 7769 9873 7803
rect 9873 7769 9907 7803
rect 9907 7769 9916 7803
rect 9864 7760 9916 7769
rect 10508 7939 10560 7948
rect 10508 7905 10517 7939
rect 10517 7905 10551 7939
rect 10551 7905 10560 7939
rect 10508 7896 10560 7905
rect 11336 7896 11388 7948
rect 11704 7896 11756 7948
rect 12624 7896 12676 7948
rect 11244 7828 11296 7880
rect 13360 7896 13412 7948
rect 10048 7735 10100 7744
rect 10048 7701 10057 7735
rect 10057 7701 10091 7735
rect 10091 7701 10100 7735
rect 10048 7692 10100 7701
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 11428 7692 11480 7744
rect 14740 7896 14792 7948
rect 15016 7939 15068 7948
rect 15016 7905 15025 7939
rect 15025 7905 15059 7939
rect 15059 7905 15068 7939
rect 15016 7896 15068 7905
rect 15108 7896 15160 7948
rect 16028 8032 16080 8084
rect 17224 8032 17276 8084
rect 21456 8075 21508 8084
rect 21456 8041 21465 8075
rect 21465 8041 21499 8075
rect 21499 8041 21508 8075
rect 21456 8032 21508 8041
rect 21824 8032 21876 8084
rect 16120 7939 16172 7948
rect 16120 7905 16129 7939
rect 16129 7905 16163 7939
rect 16163 7905 16172 7939
rect 16120 7896 16172 7905
rect 16396 7939 16448 7948
rect 16396 7905 16430 7939
rect 16430 7905 16448 7939
rect 16396 7896 16448 7905
rect 17408 7896 17460 7948
rect 17684 7939 17736 7948
rect 17684 7905 17693 7939
rect 17693 7905 17727 7939
rect 17727 7905 17736 7939
rect 17684 7896 17736 7905
rect 22652 8032 22704 8084
rect 22744 7896 22796 7948
rect 12716 7735 12768 7744
rect 12716 7701 12725 7735
rect 12725 7701 12759 7735
rect 12759 7701 12768 7735
rect 12716 7692 12768 7701
rect 12808 7692 12860 7744
rect 14832 7803 14884 7812
rect 14832 7769 14841 7803
rect 14841 7769 14875 7803
rect 14875 7769 14884 7803
rect 14832 7760 14884 7769
rect 17132 7828 17184 7880
rect 19984 7828 20036 7880
rect 15108 7760 15160 7812
rect 15844 7692 15896 7744
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 8208 7488 8260 7540
rect 8300 7488 8352 7540
rect 5816 7420 5868 7472
rect 5264 7352 5316 7404
rect 6184 7216 6236 7268
rect 8116 7420 8168 7472
rect 8944 7488 8996 7540
rect 10324 7488 10376 7540
rect 10508 7488 10560 7540
rect 11704 7531 11756 7540
rect 11704 7497 11713 7531
rect 11713 7497 11747 7531
rect 11747 7497 11756 7531
rect 11704 7488 11756 7497
rect 12532 7488 12584 7540
rect 12624 7488 12676 7540
rect 13268 7488 13320 7540
rect 14832 7488 14884 7540
rect 14924 7531 14976 7540
rect 14924 7497 14933 7531
rect 14933 7497 14967 7531
rect 14967 7497 14976 7531
rect 14924 7488 14976 7497
rect 9680 7420 9732 7472
rect 9864 7420 9916 7472
rect 9956 7463 10008 7472
rect 9956 7429 9965 7463
rect 9965 7429 9999 7463
rect 9999 7429 10008 7463
rect 9956 7420 10008 7429
rect 10048 7463 10100 7472
rect 10048 7429 10057 7463
rect 10057 7429 10091 7463
rect 10091 7429 10100 7463
rect 10048 7420 10100 7429
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 9036 7327 9088 7336
rect 7472 7216 7524 7268
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 10232 7284 10284 7336
rect 10692 7284 10744 7336
rect 11336 7284 11388 7336
rect 11428 7327 11480 7336
rect 11428 7293 11437 7327
rect 11437 7293 11471 7327
rect 11471 7293 11480 7327
rect 11428 7284 11480 7293
rect 11612 7284 11664 7336
rect 12624 7395 12676 7404
rect 12624 7361 12633 7395
rect 12633 7361 12667 7395
rect 12667 7361 12676 7395
rect 12624 7352 12676 7361
rect 14556 7420 14608 7472
rect 17408 7488 17460 7540
rect 20168 7420 20220 7472
rect 20536 7488 20588 7540
rect 22192 7488 22244 7540
rect 5632 7148 5684 7200
rect 7564 7191 7616 7200
rect 7564 7157 7573 7191
rect 7573 7157 7607 7191
rect 7607 7157 7616 7191
rect 7564 7148 7616 7157
rect 11152 7259 11204 7268
rect 11152 7225 11170 7259
rect 11170 7225 11204 7259
rect 11152 7216 11204 7225
rect 13360 7284 13412 7336
rect 14372 7284 14424 7336
rect 15844 7327 15896 7336
rect 15844 7293 15878 7327
rect 15878 7293 15896 7327
rect 12808 7148 12860 7200
rect 12992 7259 13044 7268
rect 12992 7225 13001 7259
rect 13001 7225 13035 7259
rect 13035 7225 13044 7259
rect 12992 7216 13044 7225
rect 14096 7216 14148 7268
rect 15844 7284 15896 7293
rect 16120 7284 16172 7336
rect 19524 7284 19576 7336
rect 20076 7284 20128 7336
rect 22100 7284 22152 7336
rect 22284 7284 22336 7336
rect 22836 7284 22888 7336
rect 14740 7148 14792 7200
rect 18420 7148 18472 7200
rect 19432 7148 19484 7200
rect 19800 7148 19852 7200
rect 19984 7191 20036 7200
rect 19984 7157 19993 7191
rect 19993 7157 20027 7191
rect 20027 7157 20036 7191
rect 19984 7148 20036 7157
rect 20720 7216 20772 7268
rect 22560 7216 22612 7268
rect 21640 7191 21692 7200
rect 21640 7157 21649 7191
rect 21649 7157 21683 7191
rect 21683 7157 21692 7191
rect 21640 7148 21692 7157
rect 19022 7046 19074 7098
rect 19086 7046 19138 7098
rect 19150 7046 19202 7098
rect 19214 7046 19266 7098
rect 19278 7046 19330 7098
rect 9956 6944 10008 6996
rect 10692 6944 10744 6996
rect 11152 6987 11204 6996
rect 11152 6953 11161 6987
rect 11161 6953 11195 6987
rect 11195 6953 11204 6987
rect 11152 6944 11204 6953
rect 12716 6944 12768 6996
rect 6184 6876 6236 6928
rect 7564 6876 7616 6928
rect 9680 6919 9732 6928
rect 9680 6885 9714 6919
rect 9714 6885 9732 6919
rect 9680 6876 9732 6885
rect 5908 6740 5960 6792
rect 5356 6672 5408 6724
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6552 6740 6604 6792
rect 7104 6808 7156 6860
rect 12992 6944 13044 6996
rect 14096 6987 14148 6996
rect 14096 6953 14105 6987
rect 14105 6953 14139 6987
rect 14139 6953 14148 6987
rect 14096 6944 14148 6953
rect 16396 6944 16448 6996
rect 18144 6944 18196 6996
rect 15016 6876 15068 6928
rect 15292 6876 15344 6928
rect 19708 6944 19760 6996
rect 20076 6944 20128 6996
rect 20444 6987 20496 6996
rect 20444 6953 20453 6987
rect 20453 6953 20487 6987
rect 20487 6953 20496 6987
rect 20444 6944 20496 6953
rect 20720 6944 20772 6996
rect 21364 6944 21416 6996
rect 21640 6944 21692 6996
rect 19984 6876 20036 6928
rect 20260 6919 20312 6928
rect 20260 6885 20269 6919
rect 20269 6885 20303 6919
rect 20303 6885 20312 6919
rect 20260 6876 20312 6885
rect 14004 6851 14056 6860
rect 14004 6817 14013 6851
rect 14013 6817 14047 6851
rect 14047 6817 14056 6851
rect 14004 6808 14056 6817
rect 14648 6808 14700 6860
rect 15660 6808 15712 6860
rect 4252 6604 4304 6656
rect 5172 6604 5224 6656
rect 5264 6647 5316 6656
rect 5264 6613 5273 6647
rect 5273 6613 5307 6647
rect 5307 6613 5316 6647
rect 5264 6604 5316 6613
rect 7012 6672 7064 6724
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 8576 6604 8628 6656
rect 11428 6604 11480 6656
rect 18880 6808 18932 6860
rect 19156 6808 19208 6860
rect 18788 6672 18840 6724
rect 19156 6672 19208 6724
rect 19524 6740 19576 6792
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 20352 6808 20404 6860
rect 21088 6876 21140 6928
rect 22192 6876 22244 6928
rect 22560 6987 22612 6996
rect 22560 6953 22569 6987
rect 22569 6953 22603 6987
rect 22603 6953 22612 6987
rect 22560 6944 22612 6953
rect 22744 6944 22796 6996
rect 20904 6808 20956 6860
rect 20628 6740 20680 6792
rect 19708 6672 19760 6724
rect 20812 6672 20864 6724
rect 22008 6851 22060 6860
rect 22008 6817 22017 6851
rect 22017 6817 22051 6851
rect 22051 6817 22060 6851
rect 22008 6808 22060 6817
rect 21456 6783 21508 6792
rect 21456 6749 21465 6783
rect 21465 6749 21499 6783
rect 21499 6749 21508 6783
rect 21456 6740 21508 6749
rect 21916 6740 21968 6792
rect 22468 6851 22520 6860
rect 22468 6817 22477 6851
rect 22477 6817 22511 6851
rect 22511 6817 22520 6851
rect 22468 6808 22520 6817
rect 18328 6647 18380 6656
rect 18328 6613 18337 6647
rect 18337 6613 18371 6647
rect 18371 6613 18380 6647
rect 18328 6604 18380 6613
rect 19800 6647 19852 6656
rect 19800 6613 19809 6647
rect 19809 6613 19843 6647
rect 19843 6613 19852 6647
rect 19800 6604 19852 6613
rect 20076 6604 20128 6656
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 21548 6647 21600 6656
rect 21548 6613 21557 6647
rect 21557 6613 21591 6647
rect 21591 6613 21600 6647
rect 21548 6604 21600 6613
rect 21916 6647 21968 6656
rect 21916 6613 21925 6647
rect 21925 6613 21959 6647
rect 21959 6613 21968 6647
rect 21916 6604 21968 6613
rect 22100 6604 22152 6656
rect 22744 6851 22796 6860
rect 22744 6817 22753 6851
rect 22753 6817 22787 6851
rect 22787 6817 22796 6851
rect 22744 6808 22796 6817
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 6184 6400 6236 6452
rect 6276 6400 6328 6452
rect 4344 6239 4396 6248
rect 4344 6205 4353 6239
rect 4353 6205 4387 6239
rect 4387 6205 4396 6239
rect 4344 6196 4396 6205
rect 5080 6196 5132 6248
rect 5264 6239 5316 6248
rect 5264 6205 5287 6239
rect 5287 6205 5316 6239
rect 5264 6196 5316 6205
rect 7012 6443 7064 6452
rect 7012 6409 7021 6443
rect 7021 6409 7055 6443
rect 7055 6409 7064 6443
rect 7012 6400 7064 6409
rect 18328 6400 18380 6452
rect 18880 6400 18932 6452
rect 20260 6400 20312 6452
rect 6828 6264 6880 6316
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 5908 6128 5960 6180
rect 6276 6128 6328 6180
rect 4252 6060 4304 6112
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 4896 6103 4948 6112
rect 4896 6069 4905 6103
rect 4905 6069 4939 6103
rect 4939 6069 4948 6103
rect 4896 6060 4948 6069
rect 6368 6060 6420 6112
rect 6644 6103 6696 6112
rect 6644 6069 6653 6103
rect 6653 6069 6687 6103
rect 6687 6069 6696 6103
rect 17868 6239 17920 6248
rect 17868 6205 17877 6239
rect 17877 6205 17911 6239
rect 17911 6205 17920 6239
rect 17868 6196 17920 6205
rect 19800 6332 19852 6384
rect 20536 6332 20588 6384
rect 18144 6239 18196 6248
rect 18144 6205 18153 6239
rect 18153 6205 18187 6239
rect 18187 6205 18196 6239
rect 18144 6196 18196 6205
rect 18420 6196 18472 6248
rect 18696 6239 18748 6248
rect 18696 6205 18705 6239
rect 18705 6205 18739 6239
rect 18739 6205 18748 6239
rect 18696 6196 18748 6205
rect 19892 6196 19944 6248
rect 20168 6196 20220 6248
rect 20352 6196 20404 6248
rect 21088 6307 21140 6316
rect 21088 6273 21097 6307
rect 21097 6273 21131 6307
rect 21131 6273 21140 6307
rect 21088 6264 21140 6273
rect 21456 6332 21508 6384
rect 22744 6400 22796 6452
rect 22652 6375 22704 6384
rect 22652 6341 22661 6375
rect 22661 6341 22695 6375
rect 22695 6341 22704 6375
rect 22652 6332 22704 6341
rect 22008 6264 22060 6316
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 21364 6239 21416 6248
rect 21364 6205 21373 6239
rect 21373 6205 21407 6239
rect 21407 6205 21416 6239
rect 21364 6196 21416 6205
rect 21824 6196 21876 6248
rect 21548 6128 21600 6180
rect 22100 6171 22152 6180
rect 22100 6137 22109 6171
rect 22109 6137 22143 6171
rect 22143 6137 22152 6171
rect 22100 6128 22152 6137
rect 22560 6239 22612 6248
rect 22560 6205 22569 6239
rect 22569 6205 22603 6239
rect 22603 6205 22612 6239
rect 22560 6196 22612 6205
rect 22836 6239 22888 6248
rect 22836 6205 22845 6239
rect 22845 6205 22879 6239
rect 22879 6205 22888 6239
rect 22836 6196 22888 6205
rect 6644 6060 6696 6069
rect 7380 6103 7432 6112
rect 7380 6069 7389 6103
rect 7389 6069 7423 6103
rect 7423 6069 7432 6103
rect 7380 6060 7432 6069
rect 18512 6103 18564 6112
rect 18512 6069 18521 6103
rect 18521 6069 18555 6103
rect 18555 6069 18564 6103
rect 18512 6060 18564 6069
rect 20168 6103 20220 6112
rect 20168 6069 20177 6103
rect 20177 6069 20211 6103
rect 20211 6069 20220 6103
rect 20168 6060 20220 6069
rect 21364 6060 21416 6112
rect 22008 6060 22060 6112
rect 19022 5958 19074 6010
rect 19086 5958 19138 6010
rect 19150 5958 19202 6010
rect 19214 5958 19266 6010
rect 19278 5958 19330 6010
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 4344 5856 4396 5908
rect 4896 5856 4948 5908
rect 5080 5856 5132 5908
rect 5816 5856 5868 5908
rect 6920 5856 6972 5908
rect 18512 5856 18564 5908
rect 19524 5856 19576 5908
rect 20168 5856 20220 5908
rect 20352 5856 20404 5908
rect 21824 5856 21876 5908
rect 22560 5856 22612 5908
rect 5540 5720 5592 5772
rect 5724 5720 5776 5772
rect 18696 5720 18748 5772
rect 19800 5720 19852 5772
rect 22192 5788 22244 5840
rect 21732 5763 21784 5772
rect 21732 5729 21766 5763
rect 21766 5729 21784 5763
rect 21732 5720 21784 5729
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 6828 5516 6880 5568
rect 7472 5559 7524 5568
rect 7472 5525 7481 5559
rect 7481 5525 7515 5559
rect 7515 5525 7524 5559
rect 7472 5516 7524 5525
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 5724 5312 5776 5364
rect 6368 5312 6420 5364
rect 18144 5312 18196 5364
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 21732 5312 21784 5364
rect 4528 5108 4580 5160
rect 5080 5151 5132 5160
rect 5080 5117 5089 5151
rect 5089 5117 5123 5151
rect 5123 5117 5132 5151
rect 5080 5108 5132 5117
rect 6276 5176 6328 5228
rect 6828 5176 6880 5228
rect 19800 5176 19852 5228
rect 5632 5108 5684 5160
rect 18788 5151 18840 5160
rect 18788 5117 18797 5151
rect 18797 5117 18831 5151
rect 18831 5117 18840 5151
rect 18788 5108 18840 5117
rect 18880 5108 18932 5160
rect 22008 5176 22060 5228
rect 21916 5108 21968 5160
rect 20260 5083 20312 5092
rect 20260 5049 20294 5083
rect 20294 5049 20312 5083
rect 20260 5040 20312 5049
rect 19022 4870 19074 4922
rect 19086 4870 19138 4922
rect 19150 4870 19202 4922
rect 19214 4870 19266 4922
rect 19278 4870 19330 4922
rect 5540 4768 5592 4820
rect 20260 4811 20312 4820
rect 20260 4777 20269 4811
rect 20269 4777 20303 4811
rect 20303 4777 20312 4811
rect 20260 4768 20312 4777
rect 20444 4768 20496 4820
rect 7380 4632 7432 4684
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 6644 4564 6696 4616
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 22284 4088 22336 4140
rect 23020 4063 23072 4072
rect 23020 4029 23029 4063
rect 23029 4029 23063 4063
rect 23063 4029 23072 4063
rect 23020 4020 23072 4029
rect 19022 3782 19074 3834
rect 19086 3782 19138 3834
rect 19150 3782 19202 3834
rect 19214 3782 19266 3834
rect 19278 3782 19330 3834
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 19022 2694 19074 2746
rect 19086 2694 19138 2746
rect 19150 2694 19202 2746
rect 19214 2694 19266 2746
rect 19278 2694 19330 2746
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 19022 1606 19074 1658
rect 19086 1606 19138 1658
rect 19150 1606 19202 1658
rect 19214 1606 19266 1658
rect 19278 1606 19330 1658
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 19022 518 19074 570
rect 19086 518 19138 570
rect 19150 518 19202 570
rect 19214 518 19266 570
rect 19278 518 19330 570
<< metal2 >>
rect 1674 23600 1730 24000
rect 4618 23600 4674 24000
rect 7562 23600 7618 24000
rect 10506 23600 10562 24000
rect 13450 23600 13506 24000
rect 16394 23746 16450 24000
rect 19338 23746 19394 24000
rect 16394 23718 17080 23746
rect 16394 23600 16450 23718
rect 1688 23322 1716 23600
rect 1676 23316 1728 23322
rect 1676 23258 1728 23264
rect 4632 23254 4660 23600
rect 7576 23254 7604 23600
rect 10520 23338 10548 23600
rect 10520 23310 10732 23338
rect 10704 23254 10732 23310
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 4620 23248 4672 23254
rect 4620 23190 4672 23196
rect 7564 23248 7616 23254
rect 7564 23190 7616 23196
rect 10692 23248 10744 23254
rect 10692 23190 10744 23196
rect 5816 23180 5868 23186
rect 5816 23122 5868 23128
rect 7196 23180 7248 23186
rect 7196 23122 7248 23128
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 4344 22976 4396 22982
rect 4344 22918 4396 22924
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 3662 22876 3970 22885
rect 3662 22874 3668 22876
rect 3724 22874 3748 22876
rect 3804 22874 3828 22876
rect 3884 22874 3908 22876
rect 3964 22874 3970 22876
rect 3724 22822 3726 22874
rect 3906 22822 3908 22874
rect 3662 22820 3668 22822
rect 3724 22820 3748 22822
rect 3804 22820 3828 22822
rect 3884 22820 3908 22822
rect 3964 22820 3970 22822
rect 3662 22811 3970 22820
rect 4356 22166 4384 22918
rect 4908 22574 4936 22918
rect 5828 22778 5856 23122
rect 5908 23112 5960 23118
rect 5908 23054 5960 23060
rect 5816 22772 5868 22778
rect 5816 22714 5868 22720
rect 5264 22704 5316 22710
rect 5264 22646 5316 22652
rect 4620 22568 4672 22574
rect 4620 22510 4672 22516
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 4344 22160 4396 22166
rect 4344 22102 4396 22108
rect 3662 21788 3970 21797
rect 3662 21786 3668 21788
rect 3724 21786 3748 21788
rect 3804 21786 3828 21788
rect 3884 21786 3908 21788
rect 3964 21786 3970 21788
rect 3724 21734 3726 21786
rect 3906 21734 3908 21786
rect 3662 21732 3668 21734
rect 3724 21732 3748 21734
rect 3804 21732 3828 21734
rect 3884 21732 3908 21734
rect 3964 21732 3970 21734
rect 3662 21723 3970 21732
rect 3662 20700 3970 20709
rect 3662 20698 3668 20700
rect 3724 20698 3748 20700
rect 3804 20698 3828 20700
rect 3884 20698 3908 20700
rect 3964 20698 3970 20700
rect 3724 20646 3726 20698
rect 3906 20646 3908 20698
rect 3662 20644 3668 20646
rect 3724 20644 3748 20646
rect 3804 20644 3828 20646
rect 3884 20644 3908 20646
rect 3964 20644 3970 20646
rect 3662 20635 3970 20644
rect 4356 20398 4384 22102
rect 4632 21010 4660 22510
rect 4896 22432 4948 22438
rect 4896 22374 4948 22380
rect 4908 22234 4936 22374
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 5276 22094 5304 22646
rect 5920 22574 5948 23054
rect 6644 23044 6696 23050
rect 6644 22986 6696 22992
rect 6656 22574 6684 22986
rect 7104 22976 7156 22982
rect 7104 22918 7156 22924
rect 5908 22568 5960 22574
rect 5908 22510 5960 22516
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6644 22568 6696 22574
rect 7116 22522 7144 22918
rect 7208 22710 7236 23122
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 7196 22704 7248 22710
rect 7196 22646 7248 22652
rect 6644 22510 6696 22516
rect 5920 22094 5948 22510
rect 5184 22066 5304 22094
rect 5644 22066 5948 22094
rect 6196 22094 6224 22510
rect 7024 22494 7144 22522
rect 7196 22500 7248 22506
rect 6644 22432 6696 22438
rect 6696 22392 6776 22420
rect 6644 22374 6696 22380
rect 6748 22166 6776 22392
rect 6736 22160 6788 22166
rect 6736 22102 6788 22108
rect 6196 22066 6316 22094
rect 5184 21894 5212 22066
rect 5172 21888 5224 21894
rect 5172 21830 5224 21836
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 4448 20398 4476 20878
rect 4632 20398 4660 20946
rect 5184 20806 5212 21830
rect 5356 21072 5408 21078
rect 5644 21026 5672 22066
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 5408 21020 5672 21026
rect 5356 21014 5672 21020
rect 5368 21010 5672 21014
rect 6090 21040 6146 21049
rect 5368 21004 5684 21010
rect 5368 20998 5632 21004
rect 5632 20946 5684 20952
rect 6000 21004 6052 21010
rect 6052 20984 6090 20992
rect 6052 20975 6146 20984
rect 6052 20964 6132 20975
rect 6000 20946 6052 20952
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5264 20868 5316 20874
rect 5264 20810 5316 20816
rect 5172 20800 5224 20806
rect 5172 20742 5224 20748
rect 5184 20398 5212 20742
rect 5276 20398 5304 20810
rect 5368 20398 5396 20878
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5644 20602 5672 20742
rect 5632 20596 5684 20602
rect 5632 20538 5684 20544
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 5816 20528 5868 20534
rect 5816 20470 5868 20476
rect 4344 20392 4396 20398
rect 4344 20334 4396 20340
rect 4436 20392 4488 20398
rect 4436 20334 4488 20340
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 5172 20392 5224 20398
rect 5172 20334 5224 20340
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 5356 20392 5408 20398
rect 5356 20334 5408 20340
rect 4252 20324 4304 20330
rect 4252 20266 4304 20272
rect 4264 19854 4292 20266
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 3662 19612 3970 19621
rect 3662 19610 3668 19612
rect 3724 19610 3748 19612
rect 3804 19610 3828 19612
rect 3884 19610 3908 19612
rect 3964 19610 3970 19612
rect 3724 19558 3726 19610
rect 3906 19558 3908 19610
rect 3662 19556 3668 19558
rect 3724 19556 3748 19558
rect 3804 19556 3828 19558
rect 3884 19556 3908 19558
rect 3964 19556 3970 19558
rect 3662 19547 3970 19556
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 3662 18459 3970 18468
rect 4264 18222 4292 19790
rect 4448 19310 4476 20334
rect 5184 19854 5212 20334
rect 5276 20058 5304 20334
rect 5368 20058 5396 20334
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 4908 19310 4936 19790
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 4436 19304 4488 19310
rect 4436 19246 4488 19252
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 4908 19174 4936 19246
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4724 18834 4752 19110
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4724 17678 4752 18770
rect 5276 18290 5304 19722
rect 5368 19514 5396 19994
rect 5736 19922 5764 20198
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5828 19310 5856 20470
rect 6012 19310 6040 20538
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5368 18290 5396 19110
rect 5552 18970 5580 19110
rect 5736 18970 5764 19246
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4908 17746 4936 18022
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 4540 14958 4568 15302
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 4172 13546 4200 13738
rect 4080 13530 4200 13546
rect 4068 13524 4200 13530
rect 4120 13518 4200 13524
rect 4068 13466 4120 13472
rect 4264 13410 4292 14214
rect 4436 13864 4488 13870
rect 4540 13818 4568 14894
rect 4908 14618 4936 17682
rect 5080 16040 5132 16046
rect 5170 16008 5226 16017
rect 5132 15988 5170 15994
rect 5080 15982 5170 15988
rect 5092 15966 5170 15982
rect 5170 15943 5226 15952
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 15706 5212 15846
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4488 13812 4568 13818
rect 4436 13806 4568 13812
rect 4448 13790 4568 13806
rect 4172 13382 4292 13410
rect 4172 13326 4200 13382
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4540 13190 4568 13790
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 4540 12782 4568 13126
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4264 12442 4292 12718
rect 5276 12442 5304 18226
rect 5368 13462 5396 18226
rect 5736 18222 5764 18906
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 6012 18290 6040 18702
rect 6104 18426 6132 20964
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 5828 17746 5856 18090
rect 6012 17882 6040 18226
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 6196 16590 6224 21286
rect 6288 21010 6316 22066
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6472 21894 6500 21966
rect 6828 21956 6880 21962
rect 6828 21898 6880 21904
rect 6368 21888 6420 21894
rect 6368 21830 6420 21836
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 6380 21146 6408 21830
rect 6368 21140 6420 21146
rect 6368 21082 6420 21088
rect 6276 21004 6328 21010
rect 6276 20946 6328 20952
rect 6368 21004 6420 21010
rect 6472 20992 6500 21830
rect 6840 21690 6868 21898
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6828 21412 6880 21418
rect 6828 21354 6880 21360
rect 6420 20964 6500 20992
rect 6368 20946 6420 20952
rect 6288 18834 6316 20946
rect 6380 20398 6408 20946
rect 6840 20942 6868 21354
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6380 16640 6408 20334
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6840 18834 6868 19858
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6932 19174 6960 19654
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6472 18222 6500 18566
rect 6932 18426 6960 19110
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6932 18290 6960 18362
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6460 18216 6512 18222
rect 6460 18158 6512 18164
rect 6472 17746 6500 18158
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 7024 16794 7052 22494
rect 7248 22460 7328 22488
rect 7196 22442 7248 22448
rect 7300 21962 7328 22460
rect 7288 21956 7340 21962
rect 7288 21898 7340 21904
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 7208 21486 7236 21830
rect 7300 21690 7328 21898
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7300 21146 7328 21626
rect 7392 21486 7420 22714
rect 7484 22506 7512 22918
rect 7668 22778 7696 23122
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 10324 23112 10376 23118
rect 10324 23054 10376 23060
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 7656 22772 7708 22778
rect 7656 22714 7708 22720
rect 8484 22772 8536 22778
rect 8484 22714 8536 22720
rect 7472 22500 7524 22506
rect 7472 22442 7524 22448
rect 7484 22166 7512 22442
rect 7472 22160 7524 22166
rect 7472 22102 7524 22108
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7392 21146 7420 21422
rect 7484 21350 7512 22102
rect 7668 21622 7696 22714
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 7932 22568 7984 22574
rect 7932 22510 7984 22516
rect 7840 22160 7892 22166
rect 7840 22102 7892 22108
rect 7748 22092 7800 22098
rect 7748 22034 7800 22040
rect 7760 21690 7788 22034
rect 7852 21962 7880 22102
rect 7840 21956 7892 21962
rect 7840 21898 7892 21904
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7944 21622 7972 22510
rect 8024 22500 8076 22506
rect 8024 22442 8076 22448
rect 8036 22234 8064 22442
rect 8128 22386 8156 22578
rect 8128 22358 8248 22386
rect 8024 22228 8076 22234
rect 8024 22170 8076 22176
rect 8220 21978 8248 22358
rect 8496 22030 8524 22714
rect 9508 22574 9536 22918
rect 9692 22778 9720 23054
rect 10140 23044 10192 23050
rect 10140 22986 10192 22992
rect 10152 22778 10180 22986
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 9036 22568 9088 22574
rect 9036 22510 9088 22516
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 9048 22234 9076 22510
rect 9496 22432 9548 22438
rect 9496 22374 9548 22380
rect 9036 22228 9088 22234
rect 9036 22170 9088 22176
rect 9220 22092 9272 22098
rect 9508 22080 9536 22374
rect 9272 22052 9536 22080
rect 9220 22034 9272 22040
rect 8036 21950 8248 21978
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 7656 21616 7708 21622
rect 7656 21558 7708 21564
rect 7932 21616 7984 21622
rect 7932 21558 7984 21564
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 7472 21344 7524 21350
rect 7472 21286 7524 21292
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7484 21010 7512 21286
rect 7760 21026 7788 21490
rect 8036 21418 8064 21950
rect 8116 21888 8168 21894
rect 8116 21830 8168 21836
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8024 21412 8076 21418
rect 8024 21354 8076 21360
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7576 20998 7788 21026
rect 7932 21004 7984 21010
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 7104 20324 7156 20330
rect 7104 20266 7156 20272
rect 7116 19786 7144 20266
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 7116 19310 7144 19722
rect 7300 19310 7328 20470
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 7392 17746 7420 18022
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6460 16652 6512 16658
rect 6380 16612 6460 16640
rect 6460 16594 6512 16600
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6196 16250 6224 16526
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 5908 16040 5960 16046
rect 5908 15982 5960 15988
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5460 15586 5488 15846
rect 5552 15706 5580 15914
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5460 15570 5580 15586
rect 5460 15564 5592 15570
rect 5460 15558 5540 15564
rect 5540 15506 5592 15512
rect 5644 14958 5672 15846
rect 5920 15706 5948 15982
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 6012 15366 6040 15846
rect 6104 15706 6132 15914
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6196 15570 6224 16186
rect 6472 16182 6500 16594
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 6644 16448 6696 16454
rect 6644 16390 6696 16396
rect 6460 16176 6512 16182
rect 6460 16118 6512 16124
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6380 15570 6408 16050
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5460 12238 5488 14350
rect 5736 14074 5764 14418
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 5552 11830 5580 12310
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5644 11694 5672 13466
rect 5736 11898 5764 14010
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12442 5948 12582
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 5460 10810 5488 11222
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5552 10674 5580 10950
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5644 10470 5672 11630
rect 5736 11218 5764 11834
rect 6012 11694 6040 15302
rect 6472 15162 6500 15982
rect 6564 15638 6592 16390
rect 6656 16046 6684 16390
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6734 16008 6790 16017
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6472 11694 6500 15098
rect 6656 15026 6684 15982
rect 6734 15943 6790 15952
rect 6748 15910 6776 15943
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6748 15570 6776 15846
rect 6840 15570 6868 16594
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6932 16114 6960 16390
rect 7576 16114 7604 20998
rect 7932 20946 7984 20952
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7668 20398 7696 20878
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 7760 20602 7788 20742
rect 7944 20602 7972 20946
rect 8036 20874 8064 21354
rect 8128 21010 8156 21830
rect 8220 21146 8248 21830
rect 9508 21486 9536 22052
rect 9692 21690 9720 22714
rect 10336 22710 10364 23054
rect 10324 22704 10376 22710
rect 10324 22646 10376 22652
rect 10140 22568 10192 22574
rect 10140 22510 10192 22516
rect 10152 22273 10180 22510
rect 10138 22264 10194 22273
rect 9956 22228 10008 22234
rect 10138 22199 10194 22208
rect 9956 22170 10008 22176
rect 9968 22098 9996 22170
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9496 21480 9548 21486
rect 9496 21422 9548 21428
rect 9784 21418 9812 22034
rect 10152 22030 10180 22199
rect 10336 22094 10364 22646
rect 10520 22234 10548 23122
rect 11244 22976 11296 22982
rect 11244 22918 11296 22924
rect 10508 22228 10560 22234
rect 10508 22170 10560 22176
rect 10336 22066 10548 22094
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 10520 21962 10548 22066
rect 10508 21956 10560 21962
rect 10508 21898 10560 21904
rect 10048 21616 10100 21622
rect 10232 21616 10284 21622
rect 10100 21564 10232 21570
rect 10048 21558 10284 21564
rect 10060 21542 10272 21558
rect 8760 21412 8812 21418
rect 8760 21354 8812 21360
rect 9772 21412 9824 21418
rect 9772 21354 9824 21360
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8116 21004 8168 21010
rect 8168 20964 8248 20992
rect 8116 20946 8168 20952
rect 8114 20904 8170 20913
rect 8024 20868 8076 20874
rect 8114 20839 8116 20848
rect 8024 20810 8076 20816
rect 8168 20839 8170 20848
rect 8116 20810 8168 20816
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7760 19922 7788 20538
rect 8220 20466 8248 20964
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7944 18970 7972 20334
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8404 19378 8432 20198
rect 8772 19922 8800 21354
rect 10244 21010 10272 21542
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 10428 21146 10456 21354
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 10888 21146 10916 21286
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10980 21010 11008 21354
rect 11164 21146 11192 21422
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 8760 19916 8812 19922
rect 8760 19858 8812 19864
rect 9128 19440 9180 19446
rect 9128 19382 9180 19388
rect 8392 19372 8444 19378
rect 8312 19332 8392 19360
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 7932 18964 7984 18970
rect 7932 18906 7984 18912
rect 8220 18834 8248 19246
rect 8312 18902 8340 19332
rect 8392 19314 8444 19320
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8404 18970 8432 19110
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 9140 18902 9168 19382
rect 8300 18896 8352 18902
rect 8300 18838 8352 18844
rect 9128 18896 9180 18902
rect 9128 18838 9180 18844
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7760 17338 7788 17478
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7852 16046 7880 18566
rect 8772 18426 8800 18770
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 9140 18290 9168 18838
rect 9416 18834 9444 20266
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 10060 19922 10088 19994
rect 10232 19984 10284 19990
rect 10232 19926 10284 19932
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9784 19378 9812 19790
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 10060 18970 10088 19858
rect 10244 19310 10272 19926
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11164 19378 11192 19858
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 10508 19236 10560 19242
rect 10508 19178 10560 19184
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 10520 18834 10548 19178
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 8220 17746 8248 18226
rect 9416 18222 9444 18770
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8312 17882 8340 18090
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8220 17202 8248 17682
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7300 15638 7328 15846
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6748 14906 6776 15506
rect 7668 15502 7696 15846
rect 7852 15502 7880 15982
rect 8036 15570 8064 16050
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 7208 15162 7236 15302
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 6932 14958 6960 15098
rect 7760 15094 7788 15302
rect 7748 15088 7800 15094
rect 7748 15030 7800 15036
rect 6920 14952 6972 14958
rect 6748 14878 6868 14906
rect 6920 14894 6972 14900
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6748 14618 6776 14758
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6748 14482 6776 14554
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6656 14346 6684 14418
rect 6644 14340 6696 14346
rect 6644 14282 6696 14288
rect 6748 13870 6776 14418
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6840 13394 6868 14878
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7024 14618 7052 14758
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7116 14482 7144 14758
rect 7300 14572 7512 14600
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7208 14278 7236 14418
rect 7300 14414 7328 14572
rect 7380 14482 7432 14488
rect 7484 14482 7512 14572
rect 7760 14482 7788 15030
rect 8220 14958 8248 15302
rect 8312 15162 8340 15302
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8312 14890 8340 15098
rect 8404 15026 8432 18022
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9416 17134 9444 17682
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9232 16726 9260 16934
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9232 16046 9260 16662
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 9048 14958 9076 15302
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 8300 14884 8352 14890
rect 8300 14826 8352 14832
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9416 14770 9444 17070
rect 9508 16522 9536 18566
rect 9876 17746 9904 18702
rect 10888 18290 10916 18906
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10888 17746 10916 18226
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10060 17202 10088 17478
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10796 16794 10824 16934
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 9496 16516 9548 16522
rect 9496 16458 9548 16464
rect 9508 16250 9536 16458
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 9876 15706 9904 15846
rect 10428 15706 10456 15846
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10980 15502 11008 18090
rect 11256 17746 11284 22918
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 11348 22166 11376 22510
rect 11336 22160 11388 22166
rect 11336 22102 11388 22108
rect 11440 21962 11468 22578
rect 11532 22098 11560 23258
rect 13464 23186 13492 23600
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 14372 23248 14424 23254
rect 14372 23190 14424 23196
rect 15200 23248 15252 23254
rect 15200 23190 15252 23196
rect 13452 23180 13504 23186
rect 13452 23122 13504 23128
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11520 22092 11572 22098
rect 11520 22034 11572 22040
rect 11704 22092 11756 22098
rect 11808 22094 11836 23054
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11992 22234 12020 22578
rect 14384 22574 14412 23190
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14372 22568 14424 22574
rect 14372 22510 14424 22516
rect 13912 22500 13964 22506
rect 13912 22442 13964 22448
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12900 22432 12952 22438
rect 12900 22374 12952 22380
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 11808 22066 11928 22094
rect 11704 22034 11756 22040
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 11716 21078 11744 22034
rect 11704 21072 11756 21078
rect 11704 21014 11756 21020
rect 11900 20942 11928 22066
rect 12452 21554 12480 22374
rect 12544 22137 12572 22374
rect 12530 22128 12586 22137
rect 12912 22094 12940 22374
rect 13084 22160 13136 22166
rect 13136 22120 13216 22148
rect 13084 22102 13136 22108
rect 12530 22063 12586 22072
rect 12820 22066 12940 22094
rect 12544 21554 12572 22063
rect 12820 21978 12848 22066
rect 12636 21950 12848 21978
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 11336 19984 11388 19990
rect 11336 19926 11388 19932
rect 11348 19258 11376 19926
rect 11624 19922 11652 20742
rect 11612 19916 11664 19922
rect 11612 19858 11664 19864
rect 11794 19544 11850 19553
rect 11794 19479 11850 19488
rect 11518 19408 11574 19417
rect 11808 19378 11836 19479
rect 11518 19343 11520 19352
rect 11572 19343 11574 19352
rect 11796 19372 11848 19378
rect 11520 19314 11572 19320
rect 11796 19314 11848 19320
rect 11348 19242 11468 19258
rect 11348 19236 11480 19242
rect 11348 19230 11428 19236
rect 11428 19178 11480 19184
rect 11796 18692 11848 18698
rect 11796 18634 11848 18640
rect 11808 18426 11836 18634
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11532 17202 11560 17478
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 11164 16658 11192 17002
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11440 16658 11468 16934
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11072 15502 11100 16594
rect 11164 16114 11192 16594
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11440 16046 11468 16594
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 7852 14550 7880 14758
rect 7840 14544 7892 14550
rect 7840 14486 7892 14492
rect 7380 14424 7432 14430
rect 7472 14476 7524 14482
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 14074 7236 14214
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 7392 13326 7420 14424
rect 7472 14418 7524 14424
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 8128 14346 8156 14758
rect 9140 14414 9168 14758
rect 9416 14742 9536 14770
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7484 12442 7512 12650
rect 7852 12442 7880 14214
rect 7944 13938 7972 14214
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8220 13394 8248 13874
rect 8312 13870 8340 14350
rect 9416 13870 9444 14554
rect 9508 14346 9536 14742
rect 9876 14482 9904 15302
rect 11440 15162 11468 15302
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9876 14074 9904 14418
rect 11440 14414 11468 15098
rect 11532 14958 11560 16730
rect 11716 15026 11744 16934
rect 11900 16590 11928 20878
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12176 19378 12204 20334
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 12268 18766 12296 19450
rect 12360 19174 12388 19790
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12544 19446 12572 19654
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12348 19168 12400 19174
rect 12348 19110 12400 19116
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12268 18290 12296 18566
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11992 17338 12020 17478
rect 12176 17338 12204 18158
rect 12360 18154 12388 18566
rect 12452 18222 12480 18634
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 12176 16454 12204 16934
rect 12544 16794 12572 17002
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12636 16658 12664 21950
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12728 21350 12756 21830
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12728 20874 12756 21286
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12716 20868 12768 20874
rect 12716 20810 12768 20816
rect 12820 20602 12848 20946
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12728 18290 12756 19110
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11808 14958 11836 15846
rect 12176 15094 12204 16390
rect 13004 15570 13032 20334
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13096 18630 13124 19994
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13096 18358 13124 18566
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 13188 17066 13216 22120
rect 13924 21690 13952 22442
rect 14384 22094 14412 22510
rect 14568 22438 14596 23054
rect 14924 23044 14976 23050
rect 14924 22986 14976 22992
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 14464 22094 14516 22098
rect 14384 22092 14516 22094
rect 14384 22066 14464 22092
rect 14464 22034 14516 22040
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 14292 21622 14320 21966
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 13912 21480 13964 21486
rect 13912 21422 13964 21428
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13280 17066 13308 21286
rect 13832 21162 13860 21422
rect 13740 21134 13860 21162
rect 13924 21146 13952 21422
rect 14004 21412 14056 21418
rect 14004 21354 14056 21360
rect 13912 21140 13964 21146
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 13372 20398 13400 21014
rect 13452 20868 13504 20874
rect 13452 20810 13504 20816
rect 13464 20466 13492 20810
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 13372 19922 13400 20334
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13464 19378 13492 20402
rect 13544 20324 13596 20330
rect 13544 20266 13596 20272
rect 13556 20058 13584 20266
rect 13740 20262 13768 21134
rect 13912 21082 13964 21088
rect 14016 21010 14044 21354
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14004 21004 14056 21010
rect 14004 20946 14056 20952
rect 14016 20398 14044 20946
rect 14004 20392 14056 20398
rect 14004 20334 14056 20340
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13556 17746 13584 18158
rect 13740 17882 13768 18158
rect 13832 17882 13860 19654
rect 14002 19408 14058 19417
rect 14002 19343 14004 19352
rect 14056 19343 14058 19352
rect 14096 19372 14148 19378
rect 14004 19314 14056 19320
rect 14096 19314 14148 19320
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13832 17134 13860 17818
rect 13924 17678 13952 18158
rect 14108 17678 14136 19314
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14108 17134 14136 17614
rect 14292 17542 14320 21286
rect 14476 20874 14504 22034
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14476 20398 14504 20810
rect 14568 20806 14596 22374
rect 14660 22098 14688 22918
rect 14936 22574 14964 22986
rect 14924 22568 14976 22574
rect 14924 22510 14976 22516
rect 15016 22500 15068 22506
rect 15016 22442 15068 22448
rect 15028 22166 15056 22442
rect 15016 22160 15068 22166
rect 15016 22102 15068 22108
rect 14648 22092 14700 22098
rect 14648 22034 14700 22040
rect 14660 21418 14688 22034
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14752 21554 14780 21830
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14648 21412 14700 21418
rect 14648 21354 14700 21360
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14648 21072 14700 21078
rect 14936 21049 14964 21286
rect 14648 21014 14700 21020
rect 14922 21040 14978 21049
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14568 20398 14596 20742
rect 14660 20398 14688 21014
rect 15212 21010 15240 23190
rect 15948 23186 15976 23462
rect 17052 23254 17080 23718
rect 19338 23718 19472 23746
rect 19338 23600 19394 23718
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 15936 23180 15988 23186
rect 15936 23122 15988 23128
rect 17500 23180 17552 23186
rect 17500 23122 17552 23128
rect 16304 23112 16356 23118
rect 17512 23066 17540 23122
rect 18432 23118 18460 23462
rect 19022 23420 19330 23429
rect 19022 23418 19028 23420
rect 19084 23418 19108 23420
rect 19164 23418 19188 23420
rect 19244 23418 19268 23420
rect 19324 23418 19330 23420
rect 19084 23366 19086 23418
rect 19266 23366 19268 23418
rect 19022 23364 19028 23366
rect 19084 23364 19108 23366
rect 19164 23364 19188 23366
rect 19244 23364 19268 23366
rect 19324 23364 19330 23366
rect 19022 23355 19330 23364
rect 19444 23186 19472 23718
rect 22282 23600 22338 24000
rect 20904 23316 20956 23322
rect 20904 23258 20956 23264
rect 20536 23248 20588 23254
rect 20536 23190 20588 23196
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 16304 23054 16356 23060
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 15384 22568 15436 22574
rect 15384 22510 15436 22516
rect 15568 22568 15620 22574
rect 15620 22528 15792 22556
rect 15568 22510 15620 22516
rect 15396 21010 15424 22510
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15580 21486 15608 22374
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 15764 21350 15792 22528
rect 16132 22098 16160 22918
rect 16316 22778 16344 23054
rect 17040 23044 17092 23050
rect 17040 22986 17092 22992
rect 17328 23038 17540 23066
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 16304 22772 16356 22778
rect 16304 22714 16356 22720
rect 16580 22500 16632 22506
rect 16580 22442 16632 22448
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16592 21486 16620 22442
rect 17052 22098 17080 22986
rect 17328 22574 17356 23038
rect 17776 22976 17828 22982
rect 17776 22918 17828 22924
rect 17788 22574 17816 22918
rect 18432 22642 18460 23054
rect 18708 22778 18736 23122
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 17408 22568 17460 22574
rect 17408 22510 17460 22516
rect 17776 22568 17828 22574
rect 17776 22510 17828 22516
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 17420 21894 17448 22510
rect 18604 22500 18656 22506
rect 18604 22442 18656 22448
rect 17500 22432 17552 22438
rect 17500 22374 17552 22380
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 17512 22098 17540 22374
rect 17592 22160 17644 22166
rect 17592 22102 17644 22108
rect 17500 22092 17552 22098
rect 17500 22034 17552 22040
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 16960 21622 16988 21830
rect 17144 21690 17172 21830
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16488 21412 16540 21418
rect 16488 21354 16540 21360
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 14922 20975 14978 20984
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15212 20602 15240 20946
rect 15764 20942 15792 21286
rect 16304 21140 16356 21146
rect 16304 21082 16356 21088
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 14660 19922 14688 20334
rect 15200 20324 15252 20330
rect 15200 20266 15252 20272
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 15212 19854 15240 20266
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15212 18970 15240 19790
rect 15396 19310 15424 20334
rect 16316 20262 16344 21082
rect 16500 21010 16528 21354
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 16592 20913 16620 20946
rect 16684 20942 16712 21286
rect 16672 20936 16724 20942
rect 16578 20904 16634 20913
rect 16672 20878 16724 20884
rect 17420 20874 17448 21830
rect 17604 21486 17632 22102
rect 17788 21622 17816 22374
rect 17866 22264 17922 22273
rect 18616 22234 18644 22442
rect 17866 22199 17868 22208
rect 17920 22199 17922 22208
rect 18604 22228 18656 22234
rect 17868 22170 17920 22176
rect 18604 22170 18656 22176
rect 17880 22030 17908 22170
rect 18708 22098 18736 22714
rect 19076 22574 19104 22918
rect 19352 22642 19380 23122
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19616 22976 19668 22982
rect 19616 22918 19668 22924
rect 19340 22636 19392 22642
rect 19392 22596 19472 22624
rect 19340 22578 19392 22584
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 19022 22332 19330 22341
rect 19022 22330 19028 22332
rect 19084 22330 19108 22332
rect 19164 22330 19188 22332
rect 19244 22330 19268 22332
rect 19324 22330 19330 22332
rect 19084 22278 19086 22330
rect 19266 22278 19268 22330
rect 19022 22276 19028 22278
rect 19084 22276 19108 22278
rect 19164 22276 19188 22278
rect 19244 22276 19268 22278
rect 19324 22276 19330 22278
rect 19022 22267 19330 22276
rect 18786 22128 18842 22137
rect 18696 22092 18748 22098
rect 19444 22098 19472 22596
rect 19524 22568 19576 22574
rect 19524 22510 19576 22516
rect 19536 22098 19564 22510
rect 19628 22166 19656 22918
rect 19904 22574 19932 23054
rect 20548 22930 20576 23190
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20732 23066 20760 23122
rect 20732 23038 20852 23066
rect 20548 22902 20760 22930
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19904 22438 19932 22510
rect 20732 22506 20760 22902
rect 20720 22500 20772 22506
rect 20720 22442 20772 22448
rect 19892 22432 19944 22438
rect 19892 22374 19944 22380
rect 19616 22160 19668 22166
rect 19616 22102 19668 22108
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 20536 22160 20588 22166
rect 20536 22102 20588 22108
rect 18786 22063 18788 22072
rect 18696 22034 18748 22040
rect 18840 22063 18842 22072
rect 19432 22092 19484 22098
rect 18788 22034 18840 22040
rect 19432 22034 19484 22040
rect 19524 22092 19576 22098
rect 19524 22034 19576 22040
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17776 21616 17828 21622
rect 17776 21558 17828 21564
rect 17592 21480 17644 21486
rect 17592 21422 17644 21428
rect 17880 21418 17908 21966
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 18156 21622 18184 21830
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 17868 21412 17920 21418
rect 17868 21354 17920 21360
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 16578 20839 16634 20848
rect 17408 20868 17460 20874
rect 17408 20810 17460 20816
rect 17420 20398 17448 20810
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 17512 20398 17540 20742
rect 17604 20398 17632 20946
rect 17972 20398 18000 20946
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15764 19514 15792 19858
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 16316 19310 16344 20198
rect 17236 20058 17264 20198
rect 17512 20058 17540 20334
rect 18064 20058 18092 20538
rect 18248 20398 18276 21286
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18248 20058 18276 20334
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18616 20058 18644 20198
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18708 19990 18736 21490
rect 18800 21486 18828 22034
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 19352 21418 19380 21966
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19444 21690 19472 21830
rect 19628 21706 19656 22102
rect 19708 22092 19760 22098
rect 19708 22034 19760 22040
rect 19432 21684 19484 21690
rect 19432 21626 19484 21632
rect 19536 21678 19656 21706
rect 19536 21418 19564 21678
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 19524 21412 19576 21418
rect 19524 21354 19576 21360
rect 19022 21244 19330 21253
rect 19022 21242 19028 21244
rect 19084 21242 19108 21244
rect 19164 21242 19188 21244
rect 19244 21242 19268 21244
rect 19324 21242 19330 21244
rect 19084 21190 19086 21242
rect 19266 21190 19268 21242
rect 19022 21188 19028 21190
rect 19084 21188 19108 21190
rect 19164 21188 19188 21190
rect 19244 21188 19268 21190
rect 19324 21188 19330 21190
rect 19022 21179 19330 21188
rect 19720 21078 19748 22034
rect 19996 21622 20024 22102
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 20260 22092 20312 22098
rect 20260 22034 20312 22040
rect 20180 21690 20208 22034
rect 20272 21962 20300 22034
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19800 21480 19852 21486
rect 19800 21422 19852 21428
rect 19812 21146 19840 21422
rect 19996 21146 20024 21558
rect 20272 21418 20300 21898
rect 20548 21554 20576 22102
rect 20732 22098 20760 22442
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 20824 22030 20852 23038
rect 20628 22024 20680 22030
rect 20812 22024 20864 22030
rect 20680 21972 20760 21978
rect 20628 21966 20760 21972
rect 20812 21966 20864 21972
rect 20640 21950 20760 21966
rect 20732 21894 20760 21950
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20548 21418 20576 21490
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20536 21412 20588 21418
rect 20536 21354 20588 21360
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 19708 21072 19760 21078
rect 19708 21014 19760 21020
rect 20732 20874 20760 21830
rect 20916 21554 20944 23258
rect 22296 23186 22324 23600
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21008 22642 21036 23054
rect 21548 22976 21600 22982
rect 21548 22918 21600 22924
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21008 22234 21036 22578
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 20996 22228 21048 22234
rect 20996 22170 21048 22176
rect 21100 22094 21128 22374
rect 21468 22098 21496 22578
rect 21560 22574 21588 22918
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21008 22066 21128 22094
rect 21456 22092 21508 22098
rect 21008 21690 21036 22066
rect 21456 22034 21508 22040
rect 21928 22030 21956 22578
rect 22008 22568 22060 22574
rect 22008 22510 22060 22516
rect 22192 22568 22244 22574
rect 22192 22510 22244 22516
rect 22020 22234 22048 22510
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 21916 22024 21968 22030
rect 21916 21966 21968 21972
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20916 21434 20944 21490
rect 21008 21486 21036 21626
rect 20824 21418 20944 21434
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 20812 21412 20944 21418
rect 20864 21406 20944 21412
rect 20812 21354 20864 21360
rect 21100 21010 21128 21830
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21192 21078 21220 21286
rect 21180 21072 21232 21078
rect 21180 21014 21232 21020
rect 21284 21010 21312 21626
rect 22112 21554 22140 22374
rect 22204 22234 22232 22510
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 21284 20874 21312 20946
rect 20720 20868 20772 20874
rect 20720 20810 20772 20816
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 19022 20156 19330 20165
rect 19022 20154 19028 20156
rect 19084 20154 19108 20156
rect 19164 20154 19188 20156
rect 19244 20154 19268 20156
rect 19324 20154 19330 20156
rect 19084 20102 19086 20154
rect 19266 20102 19268 20154
rect 19022 20100 19028 20102
rect 19084 20100 19108 20102
rect 19164 20100 19188 20102
rect 19244 20100 19268 20102
rect 19324 20100 19330 20102
rect 19022 20091 19330 20100
rect 18696 19984 18748 19990
rect 18696 19926 18748 19932
rect 20732 19922 20760 20810
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20824 20398 20852 20742
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 16670 19544 16726 19553
rect 16670 19479 16726 19488
rect 16684 19378 16712 19479
rect 17236 19446 17264 19790
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 18432 19378 18460 19654
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 14752 18426 14780 18770
rect 14936 18426 14964 18770
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 14924 18420 14976 18426
rect 14924 18362 14976 18368
rect 16408 18222 16436 18702
rect 16500 18358 16528 18770
rect 17328 18766 17356 19110
rect 17696 18902 17724 19246
rect 18708 19224 18736 19654
rect 19168 19446 19196 19654
rect 19996 19514 20024 19858
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 19156 19440 19208 19446
rect 19156 19382 19208 19388
rect 18788 19236 18840 19242
rect 18708 19196 18788 19224
rect 18788 19178 18840 19184
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18064 18970 18092 19110
rect 18616 18970 18644 19110
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 17684 18896 17736 18902
rect 17684 18838 17736 18844
rect 18800 18834 18828 19178
rect 18892 18850 18920 19382
rect 20548 19366 20760 19394
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19022 19068 19330 19077
rect 19022 19066 19028 19068
rect 19084 19066 19108 19068
rect 19164 19066 19188 19068
rect 19244 19066 19268 19068
rect 19324 19066 19330 19068
rect 19084 19014 19086 19066
rect 19266 19014 19268 19066
rect 19022 19012 19028 19014
rect 19084 19012 19108 19014
rect 19164 19012 19188 19014
rect 19244 19012 19268 19014
rect 19324 19012 19330 19014
rect 19022 19003 19330 19012
rect 19156 18964 19208 18970
rect 19294 18964 19346 18970
rect 19208 18924 19294 18952
rect 19156 18906 19208 18912
rect 19294 18906 19346 18912
rect 18892 18834 19196 18850
rect 18788 18828 18840 18834
rect 18892 18828 19208 18834
rect 18892 18822 19156 18828
rect 18788 18770 18840 18776
rect 19156 18770 19208 18776
rect 19294 18828 19346 18834
rect 19294 18770 19346 18776
rect 17316 18760 17368 18766
rect 19306 18714 19334 18770
rect 17316 18702 17368 18708
rect 16488 18352 16540 18358
rect 16488 18294 16540 18300
rect 17328 18222 17356 18702
rect 18708 18698 19334 18714
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 18696 18692 19334 18698
rect 18748 18686 19334 18692
rect 18696 18634 18748 18640
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18972 18624 19024 18630
rect 19156 18624 19208 18630
rect 19024 18584 19156 18612
rect 18972 18566 19024 18572
rect 19156 18566 19208 18572
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14292 17338 14320 17478
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14292 17202 14320 17274
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14568 17134 14596 18022
rect 15948 17882 15976 18158
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 16408 17678 16436 18158
rect 16856 18148 16908 18154
rect 16856 18090 16908 18096
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 13268 17060 13320 17066
rect 13268 17002 13320 17008
rect 14188 17060 14240 17066
rect 14188 17002 14240 17008
rect 13188 16590 13216 17002
rect 13280 16794 13308 17002
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12544 15144 12572 15438
rect 12452 15116 12572 15144
rect 12164 15088 12216 15094
rect 12164 15030 12216 15036
rect 12072 15020 12124 15026
rect 12452 15008 12480 15116
rect 12072 14962 12124 14968
rect 12360 14980 12480 15008
rect 12532 15020 12584 15026
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11532 14600 11560 14894
rect 11532 14572 11652 14600
rect 11624 14414 11652 14572
rect 11808 14498 11836 14894
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11716 14482 11836 14498
rect 11704 14476 11836 14482
rect 11756 14470 11836 14476
rect 11704 14418 11756 14424
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7944 12306 7972 13330
rect 8312 13326 8340 13806
rect 10060 13802 10088 14214
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 8588 13530 8616 13670
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 9784 13394 9812 13670
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 12986 8340 13126
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 8220 12170 8248 12582
rect 8404 12442 8432 13330
rect 10060 13326 10088 13738
rect 10244 13394 10272 13942
rect 10980 13802 11008 14282
rect 11440 14074 11468 14350
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 10980 13394 11008 13738
rect 11440 13394 11468 13874
rect 11716 13870 11744 14418
rect 11900 14278 11928 14758
rect 11992 14618 12020 14758
rect 12084 14618 12112 14962
rect 12360 14822 12388 14980
rect 12532 14962 12584 14968
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12544 14550 12572 14962
rect 13096 14890 13124 16526
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 13924 16046 13952 16390
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 13084 14884 13136 14890
rect 13084 14826 13136 14832
rect 12820 14618 12848 14826
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 13096 14550 13124 14826
rect 13188 14618 13216 15506
rect 13464 15162 13492 15506
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13912 15088 13964 15094
rect 13912 15030 13964 15036
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 12532 14544 12584 14550
rect 12532 14486 12584 14492
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11900 14090 11928 14214
rect 11900 14062 12020 14090
rect 12452 14074 12480 14418
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11808 13326 11836 13670
rect 11992 13394 12020 14062
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 13096 13870 13124 14486
rect 13268 14340 13320 14346
rect 13268 14282 13320 14288
rect 13280 13938 13308 14282
rect 13740 14278 13768 14758
rect 13924 14618 13952 15030
rect 14200 14958 14228 17002
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 16590 14412 16934
rect 14752 16794 14780 17138
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14660 16182 14688 16390
rect 14648 16176 14700 16182
rect 14648 16118 14700 16124
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14384 15706 14412 15982
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14568 15570 14596 15982
rect 14660 15570 14688 16118
rect 14936 15570 14964 16390
rect 15028 16114 15056 16934
rect 15120 16250 15148 17546
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16224 17338 16252 17478
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 15936 17060 15988 17066
rect 15936 17002 15988 17008
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15120 16046 15148 16186
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15672 15910 15700 16594
rect 15948 16046 15976 17002
rect 16592 16658 16620 18022
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16684 16522 16712 17274
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16592 16182 16620 16390
rect 16580 16176 16632 16182
rect 16580 16118 16632 16124
rect 16684 16046 16712 16458
rect 16776 16046 16804 16934
rect 16868 16794 16896 18090
rect 18800 17882 18828 18566
rect 19022 17980 19330 17989
rect 19022 17978 19028 17980
rect 19084 17978 19108 17980
rect 19164 17978 19188 17980
rect 19244 17978 19268 17980
rect 19324 17978 19330 17980
rect 19084 17926 19086 17978
rect 19266 17926 19268 17978
rect 19022 17924 19028 17926
rect 19084 17924 19108 17926
rect 19164 17924 19188 17926
rect 19244 17924 19268 17926
rect 19324 17924 19330 17926
rect 19022 17915 19330 17924
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 17500 17264 17552 17270
rect 17420 17212 17500 17218
rect 17420 17206 17552 17212
rect 17420 17190 17540 17206
rect 17420 17134 17448 17190
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16868 16590 16896 16730
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16960 16454 16988 17002
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17144 16658 17172 16934
rect 17420 16794 17448 17070
rect 18248 17066 18276 17478
rect 18800 17338 18828 17818
rect 19444 17814 19472 18702
rect 19340 17808 19392 17814
rect 19340 17750 19392 17756
rect 19432 17808 19484 17814
rect 19432 17750 19484 17756
rect 19064 17740 19116 17746
rect 19064 17682 19116 17688
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 18972 17604 19024 17610
rect 18972 17546 19024 17552
rect 18984 17338 19012 17546
rect 19076 17338 19104 17682
rect 19168 17542 19196 17682
rect 19352 17660 19380 17750
rect 19536 17660 19564 19110
rect 20364 18970 20392 19246
rect 20444 19168 20496 19174
rect 20548 19156 20576 19366
rect 20732 19310 20760 19366
rect 20824 19310 20852 20198
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21100 19378 21128 19654
rect 21192 19514 21220 20198
rect 21284 19922 21312 20810
rect 21916 20800 21968 20806
rect 21916 20742 21968 20748
rect 21928 20602 21956 20742
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 21928 20466 21956 20538
rect 22020 20534 22048 21286
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21468 19514 21496 20198
rect 22020 20058 22048 20470
rect 22572 20398 22600 21286
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 21548 19916 21600 19922
rect 21548 19858 21600 19864
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20496 19128 20576 19156
rect 20444 19110 20496 19116
rect 20352 18964 20404 18970
rect 20352 18906 20404 18912
rect 20444 18624 20496 18630
rect 20548 18612 20576 19128
rect 20640 18766 20668 19246
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20628 18624 20680 18630
rect 20548 18584 20628 18612
rect 20444 18566 20496 18572
rect 20628 18566 20680 18572
rect 20456 18426 20484 18566
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19352 17632 19564 17660
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 17052 16046 17080 16526
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14200 14618 14228 14894
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13740 13870 13768 14214
rect 13832 14074 13860 14214
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 15212 13938 15240 15370
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8496 12374 8524 12582
rect 9416 12434 9444 12650
rect 9416 12406 9628 12434
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5828 11150 5856 11494
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 4264 9518 4292 9862
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4356 9178 4384 9454
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 4908 8634 4936 8978
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5092 8430 5120 8570
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5184 8294 5212 8774
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 5276 7410 5304 10134
rect 5552 9382 5580 10406
rect 5644 10130 5672 10406
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5644 9654 5672 9930
rect 5736 9722 5764 11018
rect 5920 11014 5948 11494
rect 6012 11098 6040 11630
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6012 11082 6132 11098
rect 6012 11076 6144 11082
rect 6012 11070 6092 11076
rect 6092 11018 6144 11024
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 6196 10810 6224 11290
rect 7208 11014 7236 11494
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 6288 10810 6316 10950
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5552 8838 5580 9318
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5644 8634 5672 9590
rect 5736 9518 5764 9658
rect 5724 9512 5776 9518
rect 6104 9489 6132 9998
rect 6196 9518 6224 10746
rect 6564 10674 6592 10950
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6656 10266 6684 10542
rect 7208 10470 7236 10950
rect 7300 10606 7328 11290
rect 7564 11280 7616 11286
rect 7564 11222 7616 11228
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7576 10554 7604 11222
rect 7668 11218 7696 11630
rect 8220 11218 8248 12106
rect 8496 11218 8524 12310
rect 9600 12102 9628 12406
rect 9876 12374 9904 13126
rect 10336 12986 10364 13262
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 9968 12374 9996 12650
rect 10796 12442 10824 12718
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8588 11286 8616 11562
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8220 11098 8248 11154
rect 8220 11070 8524 11098
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7852 10742 7880 10950
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 8220 10674 8248 11070
rect 8496 11014 8524 11070
rect 8680 11014 8708 11494
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8404 10742 8432 10950
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8680 10674 8708 10950
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 7576 10538 7788 10554
rect 7576 10532 7800 10538
rect 7576 10526 7748 10532
rect 7748 10474 7800 10480
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6184 9512 6236 9518
rect 5724 9454 5776 9460
rect 6090 9480 6146 9489
rect 6184 9454 6236 9460
rect 6090 9415 6146 9424
rect 6104 9382 6132 9415
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5276 6662 5304 7346
rect 5368 6730 5396 8570
rect 5736 8566 5764 9318
rect 6196 9178 6224 9454
rect 6288 9450 6316 9930
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6564 9722 6592 9862
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 7012 9512 7064 9518
rect 7010 9480 7012 9489
rect 7064 9480 7066 9489
rect 6276 9444 6328 9450
rect 7010 9415 7066 9424
rect 6276 9386 6328 9392
rect 7024 9382 7052 9415
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6472 9178 6500 9318
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8566 5856 8774
rect 6196 8634 6224 9114
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6380 8634 6408 8978
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5828 7478 5856 8502
rect 6472 8430 6500 9114
rect 7760 9110 7788 10474
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 10266 8432 10406
rect 9048 10266 9076 10474
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9416 10266 9444 10406
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7748 9104 7800 9110
rect 7748 9046 7800 9052
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 7116 7954 7144 9046
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7576 8566 7604 8774
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7564 8560 7616 8566
rect 7616 8520 7696 8548
rect 7564 8502 7616 8508
rect 7300 8022 7328 8502
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 4264 6118 4292 6598
rect 5184 6338 5212 6598
rect 5184 6310 5304 6338
rect 5276 6254 5304 6310
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4264 5914 4292 6054
rect 4356 5914 4384 6190
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 4540 5166 4568 6054
rect 4908 5914 4936 6054
rect 5092 5914 5120 6190
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5092 5166 5120 5850
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5552 4826 5580 5714
rect 5644 5166 5672 7142
rect 5920 6882 5948 7890
rect 6184 7268 6236 7274
rect 6184 7210 6236 7216
rect 6196 6934 6224 7210
rect 5828 6854 5948 6882
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 5828 5914 5856 6854
rect 6196 6798 6224 6870
rect 7116 6866 7144 7890
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 5920 6186 5948 6734
rect 6196 6458 6224 6734
rect 6288 6458 6316 6734
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6196 6202 6224 6394
rect 6564 6202 6592 6734
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6196 6186 6316 6202
rect 5908 6180 5960 6186
rect 6196 6180 6328 6186
rect 6196 6174 6276 6180
rect 5908 6122 5960 6128
rect 6564 6174 6684 6202
rect 6276 6122 6328 6128
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5736 5370 5764 5714
rect 5828 5710 5856 5850
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 6288 5234 6316 6122
rect 6656 6118 6684 6174
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6380 5370 6408 6054
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 6288 4622 6316 5170
rect 6656 4622 6684 6054
rect 6840 5574 6868 6258
rect 6932 5914 6960 6598
rect 7024 6458 7052 6666
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 5234 6868 5510
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 7392 4690 7420 6054
rect 7484 5574 7512 7210
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 6934 7604 7142
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7668 6322 7696 8520
rect 7760 8294 7788 9046
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 7944 8634 7972 8774
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 8090 7788 8230
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 8128 7478 8156 8774
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8220 7546 8248 8434
rect 8312 7546 8340 8502
rect 8404 8498 8432 10066
rect 8588 8838 8616 10066
rect 9508 9994 9536 10406
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8404 8090 8432 8434
rect 8588 8430 8616 8774
rect 8772 8498 8800 9114
rect 9600 8838 9628 12038
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9692 10810 9720 11290
rect 10796 11218 10824 12378
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10980 11762 11008 12038
rect 11072 11898 11100 13262
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10784 11212 10836 11218
rect 10612 11172 10784 11200
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9876 10606 9904 11018
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 10060 10606 10088 10950
rect 10612 10742 10640 11172
rect 10784 11154 10836 11160
rect 10980 11082 11008 11698
rect 11348 11694 11376 12650
rect 11532 12374 11560 13126
rect 12912 12442 12940 13194
rect 14108 12850 14136 13670
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 13912 12776 13964 12782
rect 13832 12724 13912 12730
rect 13832 12718 13964 12724
rect 13832 12702 13952 12718
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 12348 12368 12400 12374
rect 13740 12322 13768 12378
rect 12348 12310 12400 12316
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11992 11354 12020 11494
rect 12360 11354 12388 12310
rect 13452 12300 13504 12306
rect 13648 12294 13768 12322
rect 13832 12306 13860 12702
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 13820 12300 13872 12306
rect 13648 12288 13676 12294
rect 13504 12260 13676 12288
rect 13452 12242 13504 12248
rect 13820 12242 13872 12248
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 13636 12096 13688 12102
rect 13688 12056 13860 12084
rect 13636 12038 13688 12044
rect 12452 11898 12480 12038
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 13832 11626 13860 12056
rect 13924 11898 13952 12582
rect 14384 12442 14412 12582
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14372 12096 14424 12102
rect 14568 12084 14596 13330
rect 14844 12714 14872 13670
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15120 12986 15148 13330
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15212 12782 15240 13670
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 14832 12708 14884 12714
rect 14832 12650 14884 12656
rect 15120 12102 15148 12718
rect 15304 12434 15332 12854
rect 15488 12850 15516 15846
rect 15672 15502 15700 15846
rect 16408 15706 16436 15982
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16684 15570 16712 15982
rect 18248 15978 18276 17002
rect 19022 16892 19330 16901
rect 19022 16890 19028 16892
rect 19084 16890 19108 16892
rect 19164 16890 19188 16892
rect 19244 16890 19268 16892
rect 19324 16890 19330 16892
rect 19084 16838 19086 16890
rect 19266 16838 19268 16890
rect 19022 16836 19028 16838
rect 19084 16836 19108 16838
rect 19164 16836 19188 16838
rect 19244 16836 19268 16838
rect 19324 16836 19330 16838
rect 19022 16827 19330 16836
rect 19444 16794 19472 17632
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19628 16658 19656 17818
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 19812 16658 19840 17070
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18236 15972 18288 15978
rect 18236 15914 18288 15920
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16592 14958 16620 15302
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16408 14550 16436 14894
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 13938 15884 14350
rect 16408 13938 16436 14486
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 14074 16804 14214
rect 17052 14074 17080 15438
rect 17420 14618 17448 15846
rect 18892 15706 18920 16390
rect 19022 15804 19330 15813
rect 19022 15802 19028 15804
rect 19084 15802 19108 15804
rect 19164 15802 19188 15804
rect 19244 15802 19268 15804
rect 19324 15802 19330 15804
rect 19084 15750 19086 15802
rect 19266 15750 19268 15802
rect 19022 15748 19028 15750
rect 19084 15748 19108 15750
rect 19164 15748 19188 15750
rect 19244 15748 19268 15750
rect 19324 15748 19330 15750
rect 19022 15739 19330 15748
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17788 15162 17816 15438
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 15856 12850 15884 13874
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15948 13190 15976 13670
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15304 12406 15424 12434
rect 15396 12306 15424 12406
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 14424 12056 14596 12084
rect 15108 12096 15160 12102
rect 14372 12038 14424 12044
rect 15108 12038 15160 12044
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15120 11898 15148 12038
rect 15212 11898 15240 12038
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 11520 11144 11572 11150
rect 12360 11098 12388 11290
rect 13924 11218 13952 11834
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 11520 11086 11572 11092
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10980 10810 11008 11018
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10612 10606 10640 10678
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9692 10266 9720 10474
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 10266 9812 10406
rect 10704 10266 10732 10610
rect 10980 10606 11008 10746
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8404 7342 8432 8026
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8588 6662 8616 8366
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8956 7546 8984 7890
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 9048 7342 9076 8366
rect 9600 8022 9628 8774
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10152 8498 10180 8570
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9876 7478 9904 7754
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10060 7478 10088 7686
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 10048 7472 10100 7478
rect 10152 7449 10180 8434
rect 10520 8430 10548 10066
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10612 9722 10640 9862
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 11072 9586 11100 10406
rect 11256 10266 11284 10406
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11164 9586 11192 9862
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 10048 7414 10100 7420
rect 10138 7440 10194 7449
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9692 6934 9720 7414
rect 9968 7002 9996 7414
rect 10138 7375 10194 7384
rect 10244 7342 10272 8230
rect 10520 7954 10548 8230
rect 10704 8022 10732 8298
rect 10796 8022 10824 8434
rect 10980 8430 11008 9454
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10980 8090 11008 8366
rect 11072 8294 11100 9386
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10336 7546 10364 7686
rect 10520 7546 10548 7890
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10704 7342 10732 7958
rect 11256 7886 11284 8366
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 7954 11376 8230
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11348 7342 11376 7890
rect 11428 7744 11480 7750
rect 11532 7732 11560 11086
rect 12268 11070 12388 11098
rect 12268 11014 12296 11070
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 11900 10674 11928 10950
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 12636 10606 12664 11154
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14016 10606 14044 10950
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14108 10538 14136 11154
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14200 10674 14228 10950
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14292 10606 14320 11154
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11716 9518 11744 9930
rect 12820 9586 12848 10406
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13740 8566 13768 9454
rect 13924 8974 13952 10406
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14108 9178 14136 10066
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14200 9722 14228 9862
rect 14292 9722 14320 9998
rect 14476 9722 14504 10066
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 12532 8560 12584 8566
rect 13728 8560 13780 8566
rect 12532 8502 12584 8508
rect 13634 8528 13690 8537
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11480 7704 11560 7732
rect 11428 7686 11480 7692
rect 11440 7342 11468 7686
rect 11624 7342 11652 8230
rect 12544 8090 12572 8502
rect 13728 8502 13780 8508
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 13634 8463 13636 8472
rect 13688 8463 13690 8472
rect 13636 8434 13688 8440
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12728 8090 12756 8230
rect 13188 8090 13216 8366
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13740 8090 13768 8230
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11716 7546 11744 7890
rect 12544 7546 12572 8026
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12636 7546 12664 7890
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12622 7440 12678 7449
rect 12622 7375 12624 7384
rect 12676 7375 12678 7384
rect 12624 7346 12676 7352
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 10704 7002 10732 7278
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11164 7002 11192 7210
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 11440 6662 11468 7278
rect 12728 7002 12756 7686
rect 12820 7206 12848 7686
rect 13280 7546 13308 8026
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13372 7342 13400 7890
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 13004 7002 13032 7210
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 14016 6866 14044 8502
rect 14200 8090 14228 9454
rect 14568 8906 14596 11494
rect 14752 11218 14780 11494
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 15028 11150 15056 11562
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15120 11082 15148 11834
rect 15948 11762 15976 13126
rect 16040 12986 16068 13806
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 16132 13394 16160 13738
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 13462 16252 13670
rect 17052 13530 17080 14010
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 17604 12782 17632 13126
rect 17696 12986 17724 14758
rect 18432 14618 18460 15506
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17788 14074 17816 14418
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 16316 11762 16344 12310
rect 16960 12306 16988 12718
rect 17224 12708 17276 12714
rect 17224 12650 17276 12656
rect 17236 12306 17264 12650
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 15304 11218 15332 11698
rect 16316 11354 16344 11698
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16408 11218 16436 11698
rect 16868 11694 16896 12174
rect 16960 11694 16988 12242
rect 17236 11830 17264 12242
rect 17696 12238 17724 12922
rect 17788 12782 17816 14010
rect 18432 13190 18460 14554
rect 18708 14482 18736 14894
rect 19022 14716 19330 14725
rect 19022 14714 19028 14716
rect 19084 14714 19108 14716
rect 19164 14714 19188 14716
rect 19244 14714 19268 14716
rect 19324 14714 19330 14716
rect 19084 14662 19086 14714
rect 19266 14662 19268 14714
rect 19022 14660 19028 14662
rect 19084 14660 19108 14662
rect 19164 14660 19188 14662
rect 19244 14660 19268 14662
rect 19324 14660 19330 14662
rect 19022 14651 19330 14660
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 19444 14278 19472 15438
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19616 15360 19668 15366
rect 19812 15314 19840 16594
rect 20088 15706 20116 16934
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 19616 15302 19668 15308
rect 19536 14958 19564 15302
rect 19628 15162 19656 15302
rect 19720 15286 19840 15314
rect 19616 15156 19668 15162
rect 19616 15098 19668 15104
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19444 14074 19472 14214
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19444 13954 19472 14010
rect 19352 13926 19472 13954
rect 19352 13870 19380 13926
rect 19536 13870 19564 14758
rect 19720 14482 19748 15286
rect 19996 15162 20024 15506
rect 19984 15156 20036 15162
rect 19812 15116 19984 15144
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19022 13628 19330 13637
rect 19022 13626 19028 13628
rect 19084 13626 19108 13628
rect 19164 13626 19188 13628
rect 19244 13626 19268 13628
rect 19324 13626 19330 13628
rect 19084 13574 19086 13626
rect 19266 13574 19268 13626
rect 19022 13572 19028 13574
rect 19084 13572 19108 13574
rect 19164 13572 19188 13574
rect 19244 13572 19268 13574
rect 19324 13572 19330 13574
rect 19022 13563 19330 13572
rect 19812 13462 19840 15116
rect 19984 15098 20036 15104
rect 20272 14890 20300 17682
rect 20364 17134 20392 18022
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20548 17134 20576 17614
rect 20640 17542 20668 18566
rect 20732 18358 20760 19110
rect 20720 18352 20772 18358
rect 20720 18294 20772 18300
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20732 17678 20760 18158
rect 20824 17882 20852 18158
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 21008 17746 21036 19110
rect 21100 18766 21128 19314
rect 21192 18970 21220 19450
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21376 18834 21404 19246
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21376 18154 21404 18566
rect 21456 18216 21508 18222
rect 21456 18158 21508 18164
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21376 17746 21404 18090
rect 21468 17882 21496 18158
rect 21456 17876 21508 17882
rect 21456 17818 21508 17824
rect 21560 17746 21588 19858
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 21652 18426 21680 19450
rect 22204 19242 22232 19654
rect 22296 19310 22324 20198
rect 22558 19680 22614 19689
rect 22558 19615 22614 19624
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22192 19236 22244 19242
rect 22192 19178 22244 19184
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 21836 18426 21864 19110
rect 22112 18426 22140 19110
rect 22572 18970 22600 19615
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22192 18828 22244 18834
rect 22192 18770 22244 18776
rect 22204 18442 22232 18770
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 22100 18420 22152 18426
rect 22204 18414 22416 18442
rect 22100 18362 22152 18368
rect 22112 18290 22324 18306
rect 22100 18284 22324 18290
rect 22152 18278 22324 18284
rect 22100 18226 22152 18232
rect 21824 18148 21876 18154
rect 21824 18090 21876 18096
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21732 18080 21784 18086
rect 21732 18022 21784 18028
rect 20996 17740 21048 17746
rect 20996 17682 21048 17688
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21548 17740 21600 17746
rect 21548 17682 21600 17688
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20260 14884 20312 14890
rect 20260 14826 20312 14832
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20180 14618 20208 14758
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20548 13870 20576 17070
rect 20732 14958 20760 17614
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 21100 17338 21128 17478
rect 21376 17338 21404 17546
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21192 16590 21220 17070
rect 21652 16726 21680 18022
rect 21744 17814 21772 18022
rect 21836 17882 21864 18090
rect 21824 17876 21876 17882
rect 21876 17836 21956 17864
rect 21824 17818 21876 17824
rect 21732 17808 21784 17814
rect 21732 17750 21784 17756
rect 21744 17134 21772 17750
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 21192 15638 21220 16526
rect 21928 16096 21956 17836
rect 22296 17814 22324 18278
rect 22284 17808 22336 17814
rect 22284 17750 22336 17756
rect 22388 17660 22416 18414
rect 22652 18352 22704 18358
rect 22652 18294 22704 18300
rect 22112 17632 22416 17660
rect 22112 16250 22140 17632
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 21928 16068 22140 16096
rect 22008 15972 22060 15978
rect 22008 15914 22060 15920
rect 21180 15632 21232 15638
rect 21180 15574 21232 15580
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21376 15162 21404 15506
rect 22020 15366 22048 15914
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20732 14006 20760 14894
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 14482 21496 14758
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 21456 14476 21508 14482
rect 21456 14418 21508 14424
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 21548 14408 21600 14414
rect 21652 14396 21680 14554
rect 21600 14368 21680 14396
rect 21548 14350 21600 14356
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 21008 13870 21036 14350
rect 21456 14340 21508 14346
rect 21456 14282 21508 14288
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21192 13938 21220 14214
rect 21468 14074 21496 14282
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21180 13932 21232 13938
rect 21456 13932 21508 13938
rect 21232 13892 21312 13920
rect 21180 13874 21232 13880
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 19800 13456 19852 13462
rect 19800 13398 19852 13404
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 18788 13252 18840 13258
rect 18788 13194 18840 13200
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18800 12850 18828 13194
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17788 12306 17816 12718
rect 18800 12306 18828 12786
rect 19352 12782 19380 13330
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19022 12540 19330 12549
rect 19022 12538 19028 12540
rect 19084 12538 19108 12540
rect 19164 12538 19188 12540
rect 19244 12538 19268 12540
rect 19324 12538 19330 12540
rect 19084 12486 19086 12538
rect 19266 12486 19268 12538
rect 19022 12484 19028 12486
rect 19084 12484 19108 12486
rect 19164 12484 19188 12486
rect 19244 12484 19268 12486
rect 19324 12484 19330 12486
rect 19022 12475 19330 12484
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 18788 12300 18840 12306
rect 18788 12242 18840 12248
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18248 11898 18276 12038
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 19444 11762 19472 12786
rect 20088 12434 20116 13126
rect 20364 12442 20392 13806
rect 20444 13796 20496 13802
rect 20444 13738 20496 13744
rect 20456 13394 20484 13738
rect 20548 13530 20576 13806
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20732 12986 20760 13466
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20824 12782 20852 13194
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 19904 12406 20116 12434
rect 20352 12436 20404 12442
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16224 10674 16252 10950
rect 16776 10674 16804 10950
rect 16868 10674 16896 11494
rect 16960 11354 16988 11494
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14844 9586 14872 10406
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14476 8430 14504 8774
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14384 7342 14412 8230
rect 14568 7478 14596 8842
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14646 8528 14702 8537
rect 14646 8463 14648 8472
rect 14700 8463 14702 8472
rect 14648 8434 14700 8440
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14108 7002 14136 7210
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14660 6866 14688 8298
rect 14752 7954 14780 8570
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14752 7206 14780 7890
rect 14844 7818 14872 8366
rect 14936 8294 14964 9046
rect 16040 8566 16068 10542
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16500 9178 16528 9318
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 14844 7546 14872 7754
rect 14936 7546 14964 8230
rect 15120 7954 15148 8366
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 15028 6934 15056 7890
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 15120 7698 15148 7754
rect 15304 7698 15332 8230
rect 15120 7670 15332 7698
rect 15304 6934 15332 7670
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 15292 6928 15344 6934
rect 15292 6870 15344 6876
rect 15672 6866 15700 8502
rect 16040 8362 16068 8502
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 16040 8090 16068 8298
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16132 7954 16160 8774
rect 16684 8634 16712 10542
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16868 9042 16896 9454
rect 17328 9178 17356 10542
rect 18064 10266 18092 10542
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 17866 9480 17922 9489
rect 17684 9444 17736 9450
rect 17866 9415 17922 9424
rect 17972 9450 18184 9466
rect 17972 9444 18196 9450
rect 17972 9438 18144 9444
rect 17684 9386 17736 9392
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16684 8498 16712 8570
rect 16868 8498 16896 8978
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 17236 8090 17264 8570
rect 17328 8498 17356 9114
rect 17696 8634 17724 9386
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17880 8566 17908 9415
rect 17972 9178 18000 9438
rect 18144 9386 18196 9392
rect 18248 9178 18276 9590
rect 18800 9518 18828 11562
rect 19022 11452 19330 11461
rect 19022 11450 19028 11452
rect 19084 11450 19108 11452
rect 19164 11450 19188 11452
rect 19244 11450 19268 11452
rect 19324 11450 19330 11452
rect 19084 11398 19086 11450
rect 19266 11398 19268 11450
rect 19022 11396 19028 11398
rect 19084 11396 19108 11398
rect 19164 11396 19188 11398
rect 19244 11396 19268 11398
rect 19324 11396 19330 11398
rect 19022 11387 19330 11396
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 18892 9926 18920 11154
rect 19022 10364 19330 10373
rect 19022 10362 19028 10364
rect 19084 10362 19108 10364
rect 19164 10362 19188 10364
rect 19244 10362 19268 10364
rect 19324 10362 19330 10364
rect 19084 10310 19086 10362
rect 19266 10310 19268 10362
rect 19022 10308 19028 10310
rect 19084 10308 19108 10310
rect 19164 10308 19188 10310
rect 19244 10308 19268 10310
rect 19324 10308 19330 10310
rect 19022 10299 19330 10308
rect 18880 9920 18932 9926
rect 18880 9862 18932 9868
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9586 19288 9862
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19536 9518 19564 11630
rect 19904 11218 19932 12406
rect 20732 12434 20760 12582
rect 20732 12406 20852 12434
rect 20352 12378 20404 12384
rect 20824 12306 20852 12406
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20916 11898 20944 12242
rect 21008 12238 21036 12854
rect 21192 12782 21220 13398
rect 21284 13394 21312 13892
rect 21456 13874 21508 13880
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 21100 12374 21128 12582
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 21284 12102 21312 13126
rect 21468 12986 21496 13874
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19996 11354 20024 11562
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19628 10130 19656 10950
rect 20272 10810 20300 11630
rect 20996 11552 21048 11558
rect 20996 11494 21048 11500
rect 21008 11354 21036 11494
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 21008 11098 21036 11290
rect 21376 11286 21404 12650
rect 21468 11898 21496 12718
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20548 10810 20576 11018
rect 20916 10810 20944 11086
rect 21008 11070 21128 11098
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 21008 10810 21036 10950
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 19340 9512 19392 9518
rect 19524 9512 19576 9518
rect 19392 9472 19524 9500
rect 19340 9454 19392 9460
rect 19524 9454 19576 9460
rect 18708 9178 18736 9454
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18800 9110 18828 9454
rect 19022 9276 19330 9285
rect 19022 9274 19028 9276
rect 19084 9274 19108 9276
rect 19164 9274 19188 9276
rect 19244 9274 19268 9276
rect 19324 9274 19330 9276
rect 19084 9222 19086 9274
rect 19266 9222 19268 9274
rect 19022 9220 19028 9222
rect 19084 9220 19108 9222
rect 19164 9220 19188 9222
rect 19244 9220 19268 9222
rect 19324 9220 19330 9222
rect 19022 9211 19330 9220
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 19430 9072 19486 9081
rect 19430 9007 19486 9016
rect 19444 8974 19472 9007
rect 19536 8974 19564 9454
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 8634 18092 8774
rect 18156 8634 18184 8910
rect 19628 8634 19656 10066
rect 19720 9722 19748 10066
rect 19904 9722 19932 10066
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 19708 9716 19760 9722
rect 19708 9658 19760 9664
rect 19892 9716 19944 9722
rect 19892 9658 19944 9664
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19720 9110 19748 9318
rect 19708 9104 19760 9110
rect 19708 9046 19760 9052
rect 19800 9104 19852 9110
rect 19800 9046 19852 9052
rect 19720 8974 19748 9046
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19720 8634 19748 8910
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 17868 8560 17920 8566
rect 17866 8528 17868 8537
rect 17920 8528 17922 8537
rect 17316 8492 17368 8498
rect 17866 8463 17922 8472
rect 17316 8434 17368 8440
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17420 7954 17448 8298
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17696 7954 17724 8230
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15856 7342 15884 7686
rect 16132 7342 16160 7890
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 16408 7002 16436 7890
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17144 7449 17172 7822
rect 17420 7546 17448 7890
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17130 7440 17186 7449
rect 17130 7375 17186 7384
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 17880 6254 17908 8463
rect 18708 8430 18736 8570
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18156 6254 18184 6938
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18340 6458 18368 6598
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18432 6254 18460 7142
rect 18708 6254 18736 8366
rect 19022 8188 19330 8197
rect 19022 8186 19028 8188
rect 19084 8186 19108 8188
rect 19164 8186 19188 8188
rect 19244 8186 19268 8188
rect 19324 8186 19330 8188
rect 19084 8134 19086 8186
rect 19266 8134 19268 8186
rect 19022 8132 19028 8134
rect 19084 8132 19108 8134
rect 19164 8132 19188 8134
rect 19244 8132 19268 8134
rect 19324 8132 19330 8134
rect 19022 8123 19330 8132
rect 19812 7834 19840 9046
rect 20088 9042 20116 9590
rect 20168 9512 20220 9518
rect 20166 9480 20168 9489
rect 20220 9480 20222 9489
rect 20166 9415 20222 9424
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19996 7886 20024 8842
rect 20180 8838 20208 9318
rect 20364 9042 20392 9386
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20548 8430 20576 9930
rect 20640 9926 20668 10406
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20732 9722 20760 10678
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 20916 10266 20944 10474
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20824 9602 20852 9658
rect 20732 9574 20852 9602
rect 20628 9512 20680 9518
rect 20732 9500 20760 9574
rect 20680 9472 20760 9500
rect 20628 9454 20680 9460
rect 20916 9382 20944 9998
rect 21100 9518 21128 11070
rect 21376 10470 21404 11222
rect 21468 10606 21496 11834
rect 21548 10736 21600 10742
rect 21548 10678 21600 10684
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 21376 10130 21404 10406
rect 21560 10130 21588 10678
rect 21744 10130 21772 12718
rect 21928 12442 21956 14962
rect 22020 14958 22048 15302
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 22112 14482 22140 16068
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 22112 13870 22140 14418
rect 22204 14278 22232 17206
rect 22664 16794 22692 18294
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22388 14822 22416 16050
rect 22664 14958 22692 16730
rect 23032 16658 23060 17614
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 23032 16250 23060 16594
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 22836 16040 22888 16046
rect 22836 15982 22888 15988
rect 22848 15638 22876 15982
rect 22836 15632 22888 15638
rect 22836 15574 22888 15580
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22468 14884 22520 14890
rect 22468 14826 22520 14832
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22204 14074 22232 14214
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 22112 12102 22140 12854
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 22204 12306 22232 12582
rect 22388 12434 22416 14758
rect 22480 14618 22508 14826
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22480 12850 22508 14214
rect 22664 12850 22692 14214
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 22388 12406 22508 12434
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 22296 11778 22324 12242
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22204 11750 22324 11778
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22020 10538 22048 11222
rect 22112 10606 22140 11290
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21732 10124 21784 10130
rect 21732 10066 21784 10072
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20640 8634 20668 8774
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20732 8106 20760 9318
rect 20824 8566 20852 9318
rect 20916 9178 20944 9318
rect 21100 9178 21128 9454
rect 21376 9450 21404 9862
rect 21364 9444 21416 9450
rect 21364 9386 21416 9392
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 21100 8294 21128 9114
rect 21284 9081 21312 9114
rect 21270 9072 21326 9081
rect 21270 9007 21326 9016
rect 21284 8974 21312 9007
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21560 8498 21588 10066
rect 21744 9722 21772 10066
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 21744 8498 21772 9658
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21836 8498 21864 8570
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 20732 8078 20852 8106
rect 21836 8090 21864 8434
rect 22020 8378 22048 8978
rect 21928 8350 22048 8378
rect 22112 8362 22140 9318
rect 22100 8356 22152 8362
rect 19720 7806 19840 7834
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19524 7336 19576 7342
rect 19524 7278 19576 7284
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19022 7100 19330 7109
rect 19022 7098 19028 7100
rect 19084 7098 19108 7100
rect 19164 7098 19188 7100
rect 19244 7098 19268 7100
rect 19324 7098 19330 7100
rect 19084 7046 19086 7098
rect 19266 7046 19268 7098
rect 19022 7044 19028 7046
rect 19084 7044 19108 7046
rect 19164 7044 19188 7046
rect 19244 7044 19268 7046
rect 19324 7044 19330 7046
rect 19022 7035 19330 7044
rect 19444 6914 19472 7142
rect 19260 6886 19472 6914
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 19156 6860 19208 6866
rect 19260 6848 19288 6886
rect 19208 6820 19288 6848
rect 19156 6802 19208 6808
rect 18788 6724 18840 6730
rect 18788 6666 18840 6672
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 18156 5370 18184 6190
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18524 5914 18552 6054
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18708 5778 18736 6190
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18800 5166 18828 6666
rect 18892 6458 18920 6802
rect 19168 6730 19196 6802
rect 19536 6798 19564 7278
rect 19720 7002 19748 7806
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20168 7472 20220 7478
rect 19904 7420 20168 7426
rect 19904 7414 20220 7420
rect 19904 7398 20208 7414
rect 19800 7200 19852 7206
rect 19800 7142 19852 7148
rect 19708 6996 19760 7002
rect 19708 6938 19760 6944
rect 19706 6896 19762 6905
rect 19706 6831 19762 6840
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19156 6724 19208 6730
rect 19156 6666 19208 6672
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18892 5166 18920 6394
rect 19022 6012 19330 6021
rect 19022 6010 19028 6012
rect 19084 6010 19108 6012
rect 19164 6010 19188 6012
rect 19244 6010 19268 6012
rect 19324 6010 19330 6012
rect 19084 5958 19086 6010
rect 19266 5958 19268 6010
rect 19022 5956 19028 5958
rect 19084 5956 19108 5958
rect 19164 5956 19188 5958
rect 19244 5956 19268 5958
rect 19324 5956 19330 5958
rect 19022 5947 19330 5956
rect 19536 5914 19564 6734
rect 19720 6730 19748 6831
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19812 6662 19840 7142
rect 19904 6866 19932 7398
rect 20076 7336 20128 7342
rect 20128 7296 20208 7324
rect 20076 7278 20128 7284
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19996 6934 20024 7142
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 19984 6928 20036 6934
rect 19984 6870 20036 6876
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 19812 6390 19840 6598
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 19904 6254 19932 6802
rect 20088 6662 20116 6938
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 20180 6254 20208 7296
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20260 6928 20312 6934
rect 20260 6870 20312 6876
rect 20272 6458 20300 6870
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20364 6254 20392 6802
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20180 5914 20208 6054
rect 20364 5914 20392 6190
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19812 5234 19840 5714
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18880 5160 18932 5166
rect 18880 5102 18932 5108
rect 20260 5092 20312 5098
rect 20260 5034 20312 5040
rect 19022 4924 19330 4933
rect 19022 4922 19028 4924
rect 19084 4922 19108 4924
rect 19164 4922 19188 4924
rect 19244 4922 19268 4924
rect 19324 4922 19330 4924
rect 19084 4870 19086 4922
rect 19266 4870 19268 4922
rect 19022 4868 19028 4870
rect 19084 4868 19108 4870
rect 19164 4868 19188 4870
rect 19244 4868 19268 4870
rect 19324 4868 19330 4870
rect 19022 4859 19330 4868
rect 20272 4826 20300 5034
rect 20456 4826 20484 6938
rect 20548 6390 20576 7482
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 20732 7002 20760 7210
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20640 6662 20668 6734
rect 20824 6730 20852 8078
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21364 6996 21416 7002
rect 21364 6938 21416 6944
rect 21088 6928 21140 6934
rect 20902 6896 20958 6905
rect 21088 6870 21140 6876
rect 20902 6831 20904 6840
rect 20956 6831 20958 6840
rect 20904 6802 20956 6808
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20824 6254 20852 6666
rect 21100 6322 21128 6870
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21376 6254 21404 6938
rect 21468 6798 21496 8026
rect 21640 7200 21692 7206
rect 21640 7142 21692 7148
rect 21652 7002 21680 7142
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21928 6798 21956 8350
rect 22100 8298 22152 8304
rect 22008 8288 22060 8294
rect 22008 8230 22060 8236
rect 22020 6866 22048 8230
rect 22204 7546 22232 11750
rect 22284 11620 22336 11626
rect 22284 11562 22336 11568
rect 22296 10810 22324 11562
rect 22388 11558 22416 12038
rect 22376 11552 22428 11558
rect 22376 11494 22428 11500
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22480 7426 22508 12406
rect 22560 11688 22612 11694
rect 22560 11630 22612 11636
rect 22572 9654 22600 11630
rect 22756 10198 22784 12718
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22572 9178 22600 9590
rect 22756 9178 22784 10134
rect 22560 9172 22612 9178
rect 22560 9114 22612 9120
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22112 7398 22508 7426
rect 22572 7426 22600 9114
rect 22756 8362 22784 9114
rect 22744 8356 22796 8362
rect 22744 8298 22796 8304
rect 22652 8288 22704 8294
rect 22652 8230 22704 8236
rect 22664 8090 22692 8230
rect 22652 8084 22704 8090
rect 22652 8026 22704 8032
rect 22744 7948 22796 7954
rect 22744 7890 22796 7896
rect 22572 7398 22692 7426
rect 22112 7342 22140 7398
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22192 6928 22244 6934
rect 22192 6870 22244 6876
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21468 6390 21496 6734
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 21456 6384 21508 6390
rect 21456 6326 21508 6332
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 21376 6118 21404 6190
rect 21560 6186 21588 6598
rect 21824 6248 21876 6254
rect 21824 6190 21876 6196
rect 21548 6180 21600 6186
rect 21548 6122 21600 6128
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21376 5370 21404 6054
rect 21836 5914 21864 6190
rect 21824 5908 21876 5914
rect 21824 5850 21876 5856
rect 21732 5772 21784 5778
rect 21732 5714 21784 5720
rect 21744 5370 21772 5714
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 21928 5166 21956 6598
rect 22020 6322 22048 6802
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 22112 6186 22140 6598
rect 22100 6180 22152 6186
rect 22100 6122 22152 6128
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22020 5234 22048 6054
rect 22204 5846 22232 6870
rect 22192 5840 22244 5846
rect 22192 5782 22244 5788
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 22296 4146 22324 7278
rect 22560 7268 22612 7274
rect 22560 7210 22612 7216
rect 22572 7002 22600 7210
rect 22560 6996 22612 7002
rect 22560 6938 22612 6944
rect 22468 6860 22520 6866
rect 22664 6848 22692 7398
rect 22756 7002 22784 7890
rect 22848 7342 22876 15574
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 23308 11801 23336 12242
rect 23294 11792 23350 11801
rect 23294 11727 23350 11736
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22520 6820 22692 6848
rect 22468 6802 22520 6808
rect 22664 6390 22692 6820
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22756 6458 22784 6802
rect 22744 6452 22796 6458
rect 22744 6394 22796 6400
rect 22652 6384 22704 6390
rect 22652 6326 22704 6332
rect 22848 6254 22876 7278
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22572 5914 22600 6190
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 23032 3913 23060 4014
rect 23018 3904 23074 3913
rect 19022 3836 19330 3845
rect 23018 3839 23074 3848
rect 19022 3834 19028 3836
rect 19084 3834 19108 3836
rect 19164 3834 19188 3836
rect 19244 3834 19268 3836
rect 19324 3834 19330 3836
rect 19084 3782 19086 3834
rect 19266 3782 19268 3834
rect 19022 3780 19028 3782
rect 19084 3780 19108 3782
rect 19164 3780 19188 3782
rect 19244 3780 19268 3782
rect 19324 3780 19330 3782
rect 19022 3771 19330 3780
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 19022 2748 19330 2757
rect 19022 2746 19028 2748
rect 19084 2746 19108 2748
rect 19164 2746 19188 2748
rect 19244 2746 19268 2748
rect 19324 2746 19330 2748
rect 19084 2694 19086 2746
rect 19266 2694 19268 2746
rect 19022 2692 19028 2694
rect 19084 2692 19108 2694
rect 19164 2692 19188 2694
rect 19244 2692 19268 2694
rect 19324 2692 19330 2694
rect 19022 2683 19330 2692
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 19022 1660 19330 1669
rect 19022 1658 19028 1660
rect 19084 1658 19108 1660
rect 19164 1658 19188 1660
rect 19244 1658 19268 1660
rect 19324 1658 19330 1660
rect 19084 1606 19086 1658
rect 19266 1606 19268 1658
rect 19022 1604 19028 1606
rect 19084 1604 19108 1606
rect 19164 1604 19188 1606
rect 19244 1604 19268 1606
rect 19324 1604 19330 1606
rect 19022 1595 19330 1604
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 19022 572 19330 581
rect 19022 570 19028 572
rect 19084 570 19108 572
rect 19164 570 19188 572
rect 19244 570 19268 572
rect 19324 570 19330 572
rect 19084 518 19086 570
rect 19266 518 19268 570
rect 19022 516 19028 518
rect 19084 516 19108 518
rect 19164 516 19188 518
rect 19244 516 19268 518
rect 19324 516 19330 518
rect 19022 507 19330 516
<< via2 >>
rect 3668 22874 3724 22876
rect 3748 22874 3804 22876
rect 3828 22874 3884 22876
rect 3908 22874 3964 22876
rect 3668 22822 3714 22874
rect 3714 22822 3724 22874
rect 3748 22822 3778 22874
rect 3778 22822 3790 22874
rect 3790 22822 3804 22874
rect 3828 22822 3842 22874
rect 3842 22822 3854 22874
rect 3854 22822 3884 22874
rect 3908 22822 3918 22874
rect 3918 22822 3964 22874
rect 3668 22820 3724 22822
rect 3748 22820 3804 22822
rect 3828 22820 3884 22822
rect 3908 22820 3964 22822
rect 3668 21786 3724 21788
rect 3748 21786 3804 21788
rect 3828 21786 3884 21788
rect 3908 21786 3964 21788
rect 3668 21734 3714 21786
rect 3714 21734 3724 21786
rect 3748 21734 3778 21786
rect 3778 21734 3790 21786
rect 3790 21734 3804 21786
rect 3828 21734 3842 21786
rect 3842 21734 3854 21786
rect 3854 21734 3884 21786
rect 3908 21734 3918 21786
rect 3918 21734 3964 21786
rect 3668 21732 3724 21734
rect 3748 21732 3804 21734
rect 3828 21732 3884 21734
rect 3908 21732 3964 21734
rect 3668 20698 3724 20700
rect 3748 20698 3804 20700
rect 3828 20698 3884 20700
rect 3908 20698 3964 20700
rect 3668 20646 3714 20698
rect 3714 20646 3724 20698
rect 3748 20646 3778 20698
rect 3778 20646 3790 20698
rect 3790 20646 3804 20698
rect 3828 20646 3842 20698
rect 3842 20646 3854 20698
rect 3854 20646 3884 20698
rect 3908 20646 3918 20698
rect 3918 20646 3964 20698
rect 3668 20644 3724 20646
rect 3748 20644 3804 20646
rect 3828 20644 3884 20646
rect 3908 20644 3964 20646
rect 6090 20984 6146 21040
rect 3668 19610 3724 19612
rect 3748 19610 3804 19612
rect 3828 19610 3884 19612
rect 3908 19610 3964 19612
rect 3668 19558 3714 19610
rect 3714 19558 3724 19610
rect 3748 19558 3778 19610
rect 3778 19558 3790 19610
rect 3790 19558 3804 19610
rect 3828 19558 3842 19610
rect 3842 19558 3854 19610
rect 3854 19558 3884 19610
rect 3908 19558 3918 19610
rect 3918 19558 3964 19610
rect 3668 19556 3724 19558
rect 3748 19556 3804 19558
rect 3828 19556 3884 19558
rect 3908 19556 3964 19558
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 5170 15952 5226 16008
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 6734 15952 6790 16008
rect 10138 22208 10194 22264
rect 8114 20868 8170 20904
rect 8114 20848 8116 20868
rect 8116 20848 8168 20868
rect 8168 20848 8170 20868
rect 12530 22072 12586 22128
rect 11794 19488 11850 19544
rect 11518 19372 11574 19408
rect 11518 19352 11520 19372
rect 11520 19352 11572 19372
rect 11572 19352 11574 19372
rect 14002 19372 14058 19408
rect 14002 19352 14004 19372
rect 14004 19352 14056 19372
rect 14056 19352 14058 19372
rect 14922 20984 14978 21040
rect 19028 23418 19084 23420
rect 19108 23418 19164 23420
rect 19188 23418 19244 23420
rect 19268 23418 19324 23420
rect 19028 23366 19074 23418
rect 19074 23366 19084 23418
rect 19108 23366 19138 23418
rect 19138 23366 19150 23418
rect 19150 23366 19164 23418
rect 19188 23366 19202 23418
rect 19202 23366 19214 23418
rect 19214 23366 19244 23418
rect 19268 23366 19278 23418
rect 19278 23366 19324 23418
rect 19028 23364 19084 23366
rect 19108 23364 19164 23366
rect 19188 23364 19244 23366
rect 19268 23364 19324 23366
rect 16578 20848 16634 20904
rect 17866 22228 17922 22264
rect 17866 22208 17868 22228
rect 17868 22208 17920 22228
rect 17920 22208 17922 22228
rect 19028 22330 19084 22332
rect 19108 22330 19164 22332
rect 19188 22330 19244 22332
rect 19268 22330 19324 22332
rect 19028 22278 19074 22330
rect 19074 22278 19084 22330
rect 19108 22278 19138 22330
rect 19138 22278 19150 22330
rect 19150 22278 19164 22330
rect 19188 22278 19202 22330
rect 19202 22278 19214 22330
rect 19214 22278 19244 22330
rect 19268 22278 19278 22330
rect 19278 22278 19324 22330
rect 19028 22276 19084 22278
rect 19108 22276 19164 22278
rect 19188 22276 19244 22278
rect 19268 22276 19324 22278
rect 18786 22092 18842 22128
rect 18786 22072 18788 22092
rect 18788 22072 18840 22092
rect 18840 22072 18842 22092
rect 19028 21242 19084 21244
rect 19108 21242 19164 21244
rect 19188 21242 19244 21244
rect 19268 21242 19324 21244
rect 19028 21190 19074 21242
rect 19074 21190 19084 21242
rect 19108 21190 19138 21242
rect 19138 21190 19150 21242
rect 19150 21190 19164 21242
rect 19188 21190 19202 21242
rect 19202 21190 19214 21242
rect 19214 21190 19244 21242
rect 19268 21190 19278 21242
rect 19278 21190 19324 21242
rect 19028 21188 19084 21190
rect 19108 21188 19164 21190
rect 19188 21188 19244 21190
rect 19268 21188 19324 21190
rect 19028 20154 19084 20156
rect 19108 20154 19164 20156
rect 19188 20154 19244 20156
rect 19268 20154 19324 20156
rect 19028 20102 19074 20154
rect 19074 20102 19084 20154
rect 19108 20102 19138 20154
rect 19138 20102 19150 20154
rect 19150 20102 19164 20154
rect 19188 20102 19202 20154
rect 19202 20102 19214 20154
rect 19214 20102 19244 20154
rect 19268 20102 19278 20154
rect 19278 20102 19324 20154
rect 19028 20100 19084 20102
rect 19108 20100 19164 20102
rect 19188 20100 19244 20102
rect 19268 20100 19324 20102
rect 16670 19488 16726 19544
rect 19028 19066 19084 19068
rect 19108 19066 19164 19068
rect 19188 19066 19244 19068
rect 19268 19066 19324 19068
rect 19028 19014 19074 19066
rect 19074 19014 19084 19066
rect 19108 19014 19138 19066
rect 19138 19014 19150 19066
rect 19150 19014 19164 19066
rect 19188 19014 19202 19066
rect 19202 19014 19214 19066
rect 19214 19014 19244 19066
rect 19268 19014 19278 19066
rect 19278 19014 19324 19066
rect 19028 19012 19084 19014
rect 19108 19012 19164 19014
rect 19188 19012 19244 19014
rect 19268 19012 19324 19014
rect 19028 17978 19084 17980
rect 19108 17978 19164 17980
rect 19188 17978 19244 17980
rect 19268 17978 19324 17980
rect 19028 17926 19074 17978
rect 19074 17926 19084 17978
rect 19108 17926 19138 17978
rect 19138 17926 19150 17978
rect 19150 17926 19164 17978
rect 19188 17926 19202 17978
rect 19202 17926 19214 17978
rect 19214 17926 19244 17978
rect 19268 17926 19278 17978
rect 19278 17926 19324 17978
rect 19028 17924 19084 17926
rect 19108 17924 19164 17926
rect 19188 17924 19244 17926
rect 19268 17924 19324 17926
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 6090 9424 6146 9480
rect 7010 9460 7012 9480
rect 7012 9460 7064 9480
rect 7064 9460 7066 9480
rect 7010 9424 7066 9460
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 19028 16890 19084 16892
rect 19108 16890 19164 16892
rect 19188 16890 19244 16892
rect 19268 16890 19324 16892
rect 19028 16838 19074 16890
rect 19074 16838 19084 16890
rect 19108 16838 19138 16890
rect 19138 16838 19150 16890
rect 19150 16838 19164 16890
rect 19188 16838 19202 16890
rect 19202 16838 19214 16890
rect 19214 16838 19244 16890
rect 19268 16838 19278 16890
rect 19278 16838 19324 16890
rect 19028 16836 19084 16838
rect 19108 16836 19164 16838
rect 19188 16836 19244 16838
rect 19268 16836 19324 16838
rect 19028 15802 19084 15804
rect 19108 15802 19164 15804
rect 19188 15802 19244 15804
rect 19268 15802 19324 15804
rect 19028 15750 19074 15802
rect 19074 15750 19084 15802
rect 19108 15750 19138 15802
rect 19138 15750 19150 15802
rect 19150 15750 19164 15802
rect 19188 15750 19202 15802
rect 19202 15750 19214 15802
rect 19214 15750 19244 15802
rect 19268 15750 19278 15802
rect 19278 15750 19324 15802
rect 19028 15748 19084 15750
rect 19108 15748 19164 15750
rect 19188 15748 19244 15750
rect 19268 15748 19324 15750
rect 10138 7384 10194 7440
rect 13634 8492 13690 8528
rect 13634 8472 13636 8492
rect 13636 8472 13688 8492
rect 13688 8472 13690 8492
rect 12622 7404 12678 7440
rect 12622 7384 12624 7404
rect 12624 7384 12676 7404
rect 12676 7384 12678 7404
rect 19028 14714 19084 14716
rect 19108 14714 19164 14716
rect 19188 14714 19244 14716
rect 19268 14714 19324 14716
rect 19028 14662 19074 14714
rect 19074 14662 19084 14714
rect 19108 14662 19138 14714
rect 19138 14662 19150 14714
rect 19150 14662 19164 14714
rect 19188 14662 19202 14714
rect 19202 14662 19214 14714
rect 19214 14662 19244 14714
rect 19268 14662 19278 14714
rect 19278 14662 19324 14714
rect 19028 14660 19084 14662
rect 19108 14660 19164 14662
rect 19188 14660 19244 14662
rect 19268 14660 19324 14662
rect 19028 13626 19084 13628
rect 19108 13626 19164 13628
rect 19188 13626 19244 13628
rect 19268 13626 19324 13628
rect 19028 13574 19074 13626
rect 19074 13574 19084 13626
rect 19108 13574 19138 13626
rect 19138 13574 19150 13626
rect 19150 13574 19164 13626
rect 19188 13574 19202 13626
rect 19202 13574 19214 13626
rect 19214 13574 19244 13626
rect 19268 13574 19278 13626
rect 19278 13574 19324 13626
rect 19028 13572 19084 13574
rect 19108 13572 19164 13574
rect 19188 13572 19244 13574
rect 19268 13572 19324 13574
rect 22558 19624 22614 19680
rect 19028 12538 19084 12540
rect 19108 12538 19164 12540
rect 19188 12538 19244 12540
rect 19268 12538 19324 12540
rect 19028 12486 19074 12538
rect 19074 12486 19084 12538
rect 19108 12486 19138 12538
rect 19138 12486 19150 12538
rect 19150 12486 19164 12538
rect 19188 12486 19202 12538
rect 19202 12486 19214 12538
rect 19214 12486 19244 12538
rect 19268 12486 19278 12538
rect 19278 12486 19324 12538
rect 19028 12484 19084 12486
rect 19108 12484 19164 12486
rect 19188 12484 19244 12486
rect 19268 12484 19324 12486
rect 14646 8492 14702 8528
rect 14646 8472 14648 8492
rect 14648 8472 14700 8492
rect 14700 8472 14702 8492
rect 17866 9424 17922 9480
rect 19028 11450 19084 11452
rect 19108 11450 19164 11452
rect 19188 11450 19244 11452
rect 19268 11450 19324 11452
rect 19028 11398 19074 11450
rect 19074 11398 19084 11450
rect 19108 11398 19138 11450
rect 19138 11398 19150 11450
rect 19150 11398 19164 11450
rect 19188 11398 19202 11450
rect 19202 11398 19214 11450
rect 19214 11398 19244 11450
rect 19268 11398 19278 11450
rect 19278 11398 19324 11450
rect 19028 11396 19084 11398
rect 19108 11396 19164 11398
rect 19188 11396 19244 11398
rect 19268 11396 19324 11398
rect 19028 10362 19084 10364
rect 19108 10362 19164 10364
rect 19188 10362 19244 10364
rect 19268 10362 19324 10364
rect 19028 10310 19074 10362
rect 19074 10310 19084 10362
rect 19108 10310 19138 10362
rect 19138 10310 19150 10362
rect 19150 10310 19164 10362
rect 19188 10310 19202 10362
rect 19202 10310 19214 10362
rect 19214 10310 19244 10362
rect 19268 10310 19278 10362
rect 19278 10310 19324 10362
rect 19028 10308 19084 10310
rect 19108 10308 19164 10310
rect 19188 10308 19244 10310
rect 19268 10308 19324 10310
rect 19028 9274 19084 9276
rect 19108 9274 19164 9276
rect 19188 9274 19244 9276
rect 19268 9274 19324 9276
rect 19028 9222 19074 9274
rect 19074 9222 19084 9274
rect 19108 9222 19138 9274
rect 19138 9222 19150 9274
rect 19150 9222 19164 9274
rect 19188 9222 19202 9274
rect 19202 9222 19214 9274
rect 19214 9222 19244 9274
rect 19268 9222 19278 9274
rect 19278 9222 19324 9274
rect 19028 9220 19084 9222
rect 19108 9220 19164 9222
rect 19188 9220 19244 9222
rect 19268 9220 19324 9222
rect 19430 9016 19486 9072
rect 17866 8508 17868 8528
rect 17868 8508 17920 8528
rect 17920 8508 17922 8528
rect 17866 8472 17922 8508
rect 17130 7384 17186 7440
rect 19028 8186 19084 8188
rect 19108 8186 19164 8188
rect 19188 8186 19244 8188
rect 19268 8186 19324 8188
rect 19028 8134 19074 8186
rect 19074 8134 19084 8186
rect 19108 8134 19138 8186
rect 19138 8134 19150 8186
rect 19150 8134 19164 8186
rect 19188 8134 19202 8186
rect 19202 8134 19214 8186
rect 19214 8134 19244 8186
rect 19268 8134 19278 8186
rect 19278 8134 19324 8186
rect 19028 8132 19084 8134
rect 19108 8132 19164 8134
rect 19188 8132 19244 8134
rect 19268 8132 19324 8134
rect 20166 9460 20168 9480
rect 20168 9460 20220 9480
rect 20220 9460 20222 9480
rect 20166 9424 20222 9460
rect 21270 9016 21326 9072
rect 19028 7098 19084 7100
rect 19108 7098 19164 7100
rect 19188 7098 19244 7100
rect 19268 7098 19324 7100
rect 19028 7046 19074 7098
rect 19074 7046 19084 7098
rect 19108 7046 19138 7098
rect 19138 7046 19150 7098
rect 19150 7046 19164 7098
rect 19188 7046 19202 7098
rect 19202 7046 19214 7098
rect 19214 7046 19244 7098
rect 19268 7046 19278 7098
rect 19278 7046 19324 7098
rect 19028 7044 19084 7046
rect 19108 7044 19164 7046
rect 19188 7044 19244 7046
rect 19268 7044 19324 7046
rect 19706 6840 19762 6896
rect 19028 6010 19084 6012
rect 19108 6010 19164 6012
rect 19188 6010 19244 6012
rect 19268 6010 19324 6012
rect 19028 5958 19074 6010
rect 19074 5958 19084 6010
rect 19108 5958 19138 6010
rect 19138 5958 19150 6010
rect 19150 5958 19164 6010
rect 19188 5958 19202 6010
rect 19202 5958 19214 6010
rect 19214 5958 19244 6010
rect 19268 5958 19278 6010
rect 19278 5958 19324 6010
rect 19028 5956 19084 5958
rect 19108 5956 19164 5958
rect 19188 5956 19244 5958
rect 19268 5956 19324 5958
rect 19028 4922 19084 4924
rect 19108 4922 19164 4924
rect 19188 4922 19244 4924
rect 19268 4922 19324 4924
rect 19028 4870 19074 4922
rect 19074 4870 19084 4922
rect 19108 4870 19138 4922
rect 19138 4870 19150 4922
rect 19150 4870 19164 4922
rect 19188 4870 19202 4922
rect 19202 4870 19214 4922
rect 19214 4870 19244 4922
rect 19268 4870 19278 4922
rect 19278 4870 19324 4922
rect 19028 4868 19084 4870
rect 19108 4868 19164 4870
rect 19188 4868 19244 4870
rect 19268 4868 19324 4870
rect 20902 6860 20958 6896
rect 20902 6840 20904 6860
rect 20904 6840 20956 6860
rect 20956 6840 20958 6860
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 23294 11736 23350 11792
rect 23018 3848 23074 3904
rect 19028 3834 19084 3836
rect 19108 3834 19164 3836
rect 19188 3834 19244 3836
rect 19268 3834 19324 3836
rect 19028 3782 19074 3834
rect 19074 3782 19084 3834
rect 19108 3782 19138 3834
rect 19138 3782 19150 3834
rect 19150 3782 19164 3834
rect 19188 3782 19202 3834
rect 19202 3782 19214 3834
rect 19214 3782 19244 3834
rect 19268 3782 19278 3834
rect 19278 3782 19324 3834
rect 19028 3780 19084 3782
rect 19108 3780 19164 3782
rect 19188 3780 19244 3782
rect 19268 3780 19324 3782
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 19028 2746 19084 2748
rect 19108 2746 19164 2748
rect 19188 2746 19244 2748
rect 19268 2746 19324 2748
rect 19028 2694 19074 2746
rect 19074 2694 19084 2746
rect 19108 2694 19138 2746
rect 19138 2694 19150 2746
rect 19150 2694 19164 2746
rect 19188 2694 19202 2746
rect 19202 2694 19214 2746
rect 19214 2694 19244 2746
rect 19268 2694 19278 2746
rect 19278 2694 19324 2746
rect 19028 2692 19084 2694
rect 19108 2692 19164 2694
rect 19188 2692 19244 2694
rect 19268 2692 19324 2694
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 19028 1658 19084 1660
rect 19108 1658 19164 1660
rect 19188 1658 19244 1660
rect 19268 1658 19324 1660
rect 19028 1606 19074 1658
rect 19074 1606 19084 1658
rect 19108 1606 19138 1658
rect 19138 1606 19150 1658
rect 19150 1606 19164 1658
rect 19188 1606 19202 1658
rect 19202 1606 19214 1658
rect 19214 1606 19244 1658
rect 19268 1606 19278 1658
rect 19278 1606 19324 1658
rect 19028 1604 19084 1606
rect 19108 1604 19164 1606
rect 19188 1604 19244 1606
rect 19268 1604 19324 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 19028 570 19084 572
rect 19108 570 19164 572
rect 19188 570 19244 572
rect 19268 570 19324 572
rect 19028 518 19074 570
rect 19074 518 19084 570
rect 19108 518 19138 570
rect 19138 518 19150 570
rect 19150 518 19164 570
rect 19188 518 19202 570
rect 19202 518 19214 570
rect 19214 518 19244 570
rect 19268 518 19278 570
rect 19278 518 19324 570
rect 19028 516 19084 518
rect 19108 516 19164 518
rect 19188 516 19244 518
rect 19268 516 19324 518
<< metal3 >>
rect 19018 23424 19334 23425
rect 19018 23360 19024 23424
rect 19088 23360 19104 23424
rect 19168 23360 19184 23424
rect 19248 23360 19264 23424
rect 19328 23360 19334 23424
rect 19018 23359 19334 23360
rect 3658 22880 3974 22881
rect 3658 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3974 22880
rect 3658 22815 3974 22816
rect 19018 22336 19334 22337
rect 19018 22272 19024 22336
rect 19088 22272 19104 22336
rect 19168 22272 19184 22336
rect 19248 22272 19264 22336
rect 19328 22272 19334 22336
rect 19018 22271 19334 22272
rect 10133 22266 10199 22269
rect 17861 22266 17927 22269
rect 10133 22264 17927 22266
rect 10133 22208 10138 22264
rect 10194 22208 17866 22264
rect 17922 22208 17927 22264
rect 10133 22206 17927 22208
rect 10133 22203 10199 22206
rect 17861 22203 17927 22206
rect 12525 22130 12591 22133
rect 18781 22130 18847 22133
rect 12525 22128 18847 22130
rect 12525 22072 12530 22128
rect 12586 22072 18786 22128
rect 18842 22072 18847 22128
rect 12525 22070 18847 22072
rect 12525 22067 12591 22070
rect 18781 22067 18847 22070
rect 3658 21792 3974 21793
rect 3658 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3974 21792
rect 3658 21727 3974 21728
rect 19018 21248 19334 21249
rect 19018 21184 19024 21248
rect 19088 21184 19104 21248
rect 19168 21184 19184 21248
rect 19248 21184 19264 21248
rect 19328 21184 19334 21248
rect 19018 21183 19334 21184
rect 6085 21042 6151 21045
rect 14917 21042 14983 21045
rect 6085 21040 14983 21042
rect 6085 20984 6090 21040
rect 6146 20984 14922 21040
rect 14978 20984 14983 21040
rect 6085 20982 14983 20984
rect 6085 20979 6151 20982
rect 14917 20979 14983 20982
rect 8109 20906 8175 20909
rect 16573 20906 16639 20909
rect 8109 20904 16639 20906
rect 8109 20848 8114 20904
rect 8170 20848 16578 20904
rect 16634 20848 16639 20904
rect 8109 20846 16639 20848
rect 8109 20843 8175 20846
rect 16573 20843 16639 20846
rect 3658 20704 3974 20705
rect 3658 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3974 20704
rect 3658 20639 3974 20640
rect 19018 20160 19334 20161
rect 19018 20096 19024 20160
rect 19088 20096 19104 20160
rect 19168 20096 19184 20160
rect 19248 20096 19264 20160
rect 19328 20096 19334 20160
rect 19018 20095 19334 20096
rect 22553 19682 22619 19685
rect 23600 19682 24000 19712
rect 22553 19680 24000 19682
rect 22553 19624 22558 19680
rect 22614 19624 24000 19680
rect 22553 19622 24000 19624
rect 22553 19619 22619 19622
rect 3658 19616 3974 19617
rect 3658 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3974 19616
rect 23600 19592 24000 19622
rect 3658 19551 3974 19552
rect 11789 19546 11855 19549
rect 16665 19546 16731 19549
rect 11789 19544 16731 19546
rect 11789 19488 11794 19544
rect 11850 19488 16670 19544
rect 16726 19488 16731 19544
rect 11789 19486 16731 19488
rect 11789 19483 11855 19486
rect 16665 19483 16731 19486
rect 11513 19410 11579 19413
rect 13997 19410 14063 19413
rect 11513 19408 14063 19410
rect 11513 19352 11518 19408
rect 11574 19352 14002 19408
rect 14058 19352 14063 19408
rect 11513 19350 14063 19352
rect 11513 19347 11579 19350
rect 13997 19347 14063 19350
rect 19018 19072 19334 19073
rect 19018 19008 19024 19072
rect 19088 19008 19104 19072
rect 19168 19008 19184 19072
rect 19248 19008 19264 19072
rect 19328 19008 19334 19072
rect 19018 19007 19334 19008
rect 3658 18528 3974 18529
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 19018 17984 19334 17985
rect 19018 17920 19024 17984
rect 19088 17920 19104 17984
rect 19168 17920 19184 17984
rect 19248 17920 19264 17984
rect 19328 17920 19334 17984
rect 19018 17919 19334 17920
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 19018 16896 19334 16897
rect 19018 16832 19024 16896
rect 19088 16832 19104 16896
rect 19168 16832 19184 16896
rect 19248 16832 19264 16896
rect 19328 16832 19334 16896
rect 19018 16831 19334 16832
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 5165 16010 5231 16013
rect 6729 16010 6795 16013
rect 5165 16008 6795 16010
rect 5165 15952 5170 16008
rect 5226 15952 6734 16008
rect 6790 15952 6795 16008
rect 5165 15950 6795 15952
rect 5165 15947 5231 15950
rect 6729 15947 6795 15950
rect 19018 15808 19334 15809
rect 19018 15744 19024 15808
rect 19088 15744 19104 15808
rect 19168 15744 19184 15808
rect 19248 15744 19264 15808
rect 19328 15744 19334 15808
rect 19018 15743 19334 15744
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 19018 14720 19334 14721
rect 19018 14656 19024 14720
rect 19088 14656 19104 14720
rect 19168 14656 19184 14720
rect 19248 14656 19264 14720
rect 19328 14656 19334 14720
rect 19018 14655 19334 14656
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 19018 13632 19334 13633
rect 19018 13568 19024 13632
rect 19088 13568 19104 13632
rect 19168 13568 19184 13632
rect 19248 13568 19264 13632
rect 19328 13568 19334 13632
rect 19018 13567 19334 13568
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 19018 12544 19334 12545
rect 19018 12480 19024 12544
rect 19088 12480 19104 12544
rect 19168 12480 19184 12544
rect 19248 12480 19264 12544
rect 19328 12480 19334 12544
rect 19018 12479 19334 12480
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 23289 11794 23355 11797
rect 23600 11794 24000 11824
rect 23289 11792 24000 11794
rect 23289 11736 23294 11792
rect 23350 11736 24000 11792
rect 23289 11734 24000 11736
rect 23289 11731 23355 11734
rect 23600 11704 24000 11734
rect 19018 11456 19334 11457
rect 19018 11392 19024 11456
rect 19088 11392 19104 11456
rect 19168 11392 19184 11456
rect 19248 11392 19264 11456
rect 19328 11392 19334 11456
rect 19018 11391 19334 11392
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 19018 10368 19334 10369
rect 19018 10304 19024 10368
rect 19088 10304 19104 10368
rect 19168 10304 19184 10368
rect 19248 10304 19264 10368
rect 19328 10304 19334 10368
rect 19018 10303 19334 10304
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 6085 9482 6151 9485
rect 7005 9482 7071 9485
rect 6085 9480 7071 9482
rect 6085 9424 6090 9480
rect 6146 9424 7010 9480
rect 7066 9424 7071 9480
rect 6085 9422 7071 9424
rect 6085 9419 6151 9422
rect 7005 9419 7071 9422
rect 17861 9482 17927 9485
rect 20161 9482 20227 9485
rect 17861 9480 20227 9482
rect 17861 9424 17866 9480
rect 17922 9424 20166 9480
rect 20222 9424 20227 9480
rect 17861 9422 20227 9424
rect 17861 9419 17927 9422
rect 20161 9419 20227 9422
rect 19018 9280 19334 9281
rect 19018 9216 19024 9280
rect 19088 9216 19104 9280
rect 19168 9216 19184 9280
rect 19248 9216 19264 9280
rect 19328 9216 19334 9280
rect 19018 9215 19334 9216
rect 19425 9074 19491 9077
rect 21265 9074 21331 9077
rect 19425 9072 21331 9074
rect 19425 9016 19430 9072
rect 19486 9016 21270 9072
rect 21326 9016 21331 9072
rect 19425 9014 21331 9016
rect 19425 9011 19491 9014
rect 21265 9011 21331 9014
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 13629 8530 13695 8533
rect 14641 8530 14707 8533
rect 17861 8530 17927 8533
rect 13629 8528 17927 8530
rect 13629 8472 13634 8528
rect 13690 8472 14646 8528
rect 14702 8472 17866 8528
rect 17922 8472 17927 8528
rect 13629 8470 17927 8472
rect 13629 8467 13695 8470
rect 14641 8467 14707 8470
rect 17861 8467 17927 8470
rect 19018 8192 19334 8193
rect 19018 8128 19024 8192
rect 19088 8128 19104 8192
rect 19168 8128 19184 8192
rect 19248 8128 19264 8192
rect 19328 8128 19334 8192
rect 19018 8127 19334 8128
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 10133 7442 10199 7445
rect 12617 7442 12683 7445
rect 17125 7442 17191 7445
rect 10133 7440 17191 7442
rect 10133 7384 10138 7440
rect 10194 7384 12622 7440
rect 12678 7384 17130 7440
rect 17186 7384 17191 7440
rect 10133 7382 17191 7384
rect 10133 7379 10199 7382
rect 12617 7379 12683 7382
rect 17125 7379 17191 7382
rect 19018 7104 19334 7105
rect 19018 7040 19024 7104
rect 19088 7040 19104 7104
rect 19168 7040 19184 7104
rect 19248 7040 19264 7104
rect 19328 7040 19334 7104
rect 19018 7039 19334 7040
rect 19701 6898 19767 6901
rect 20897 6898 20963 6901
rect 19701 6896 20963 6898
rect 19701 6840 19706 6896
rect 19762 6840 20902 6896
rect 20958 6840 20963 6896
rect 19701 6838 20963 6840
rect 19701 6835 19767 6838
rect 20897 6835 20963 6838
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 19018 6016 19334 6017
rect 19018 5952 19024 6016
rect 19088 5952 19104 6016
rect 19168 5952 19184 6016
rect 19248 5952 19264 6016
rect 19328 5952 19334 6016
rect 19018 5951 19334 5952
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 19018 4928 19334 4929
rect 19018 4864 19024 4928
rect 19088 4864 19104 4928
rect 19168 4864 19184 4928
rect 19248 4864 19264 4928
rect 19328 4864 19334 4928
rect 19018 4863 19334 4864
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 23013 3906 23079 3909
rect 23600 3906 24000 3936
rect 23013 3904 24000 3906
rect 23013 3848 23018 3904
rect 23074 3848 24000 3904
rect 23013 3846 24000 3848
rect 23013 3843 23079 3846
rect 19018 3840 19334 3841
rect 19018 3776 19024 3840
rect 19088 3776 19104 3840
rect 19168 3776 19184 3840
rect 19248 3776 19264 3840
rect 19328 3776 19334 3840
rect 23600 3816 24000 3846
rect 19018 3775 19334 3776
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 19018 2752 19334 2753
rect 19018 2688 19024 2752
rect 19088 2688 19104 2752
rect 19168 2688 19184 2752
rect 19248 2688 19264 2752
rect 19328 2688 19334 2752
rect 19018 2687 19334 2688
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 19018 1664 19334 1665
rect 19018 1600 19024 1664
rect 19088 1600 19104 1664
rect 19168 1600 19184 1664
rect 19248 1600 19264 1664
rect 19328 1600 19334 1664
rect 19018 1599 19334 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 19018 576 19334 577
rect 19018 512 19024 576
rect 19088 512 19104 576
rect 19168 512 19184 576
rect 19248 512 19264 576
rect 19328 512 19334 576
rect 19018 511 19334 512
<< via3 >>
rect 19024 23420 19088 23424
rect 19024 23364 19028 23420
rect 19028 23364 19084 23420
rect 19084 23364 19088 23420
rect 19024 23360 19088 23364
rect 19104 23420 19168 23424
rect 19104 23364 19108 23420
rect 19108 23364 19164 23420
rect 19164 23364 19168 23420
rect 19104 23360 19168 23364
rect 19184 23420 19248 23424
rect 19184 23364 19188 23420
rect 19188 23364 19244 23420
rect 19244 23364 19248 23420
rect 19184 23360 19248 23364
rect 19264 23420 19328 23424
rect 19264 23364 19268 23420
rect 19268 23364 19324 23420
rect 19324 23364 19328 23420
rect 19264 23360 19328 23364
rect 3664 22876 3728 22880
rect 3664 22820 3668 22876
rect 3668 22820 3724 22876
rect 3724 22820 3728 22876
rect 3664 22816 3728 22820
rect 3744 22876 3808 22880
rect 3744 22820 3748 22876
rect 3748 22820 3804 22876
rect 3804 22820 3808 22876
rect 3744 22816 3808 22820
rect 3824 22876 3888 22880
rect 3824 22820 3828 22876
rect 3828 22820 3884 22876
rect 3884 22820 3888 22876
rect 3824 22816 3888 22820
rect 3904 22876 3968 22880
rect 3904 22820 3908 22876
rect 3908 22820 3964 22876
rect 3964 22820 3968 22876
rect 3904 22816 3968 22820
rect 19024 22332 19088 22336
rect 19024 22276 19028 22332
rect 19028 22276 19084 22332
rect 19084 22276 19088 22332
rect 19024 22272 19088 22276
rect 19104 22332 19168 22336
rect 19104 22276 19108 22332
rect 19108 22276 19164 22332
rect 19164 22276 19168 22332
rect 19104 22272 19168 22276
rect 19184 22332 19248 22336
rect 19184 22276 19188 22332
rect 19188 22276 19244 22332
rect 19244 22276 19248 22332
rect 19184 22272 19248 22276
rect 19264 22332 19328 22336
rect 19264 22276 19268 22332
rect 19268 22276 19324 22332
rect 19324 22276 19328 22332
rect 19264 22272 19328 22276
rect 3664 21788 3728 21792
rect 3664 21732 3668 21788
rect 3668 21732 3724 21788
rect 3724 21732 3728 21788
rect 3664 21728 3728 21732
rect 3744 21788 3808 21792
rect 3744 21732 3748 21788
rect 3748 21732 3804 21788
rect 3804 21732 3808 21788
rect 3744 21728 3808 21732
rect 3824 21788 3888 21792
rect 3824 21732 3828 21788
rect 3828 21732 3884 21788
rect 3884 21732 3888 21788
rect 3824 21728 3888 21732
rect 3904 21788 3968 21792
rect 3904 21732 3908 21788
rect 3908 21732 3964 21788
rect 3964 21732 3968 21788
rect 3904 21728 3968 21732
rect 19024 21244 19088 21248
rect 19024 21188 19028 21244
rect 19028 21188 19084 21244
rect 19084 21188 19088 21244
rect 19024 21184 19088 21188
rect 19104 21244 19168 21248
rect 19104 21188 19108 21244
rect 19108 21188 19164 21244
rect 19164 21188 19168 21244
rect 19104 21184 19168 21188
rect 19184 21244 19248 21248
rect 19184 21188 19188 21244
rect 19188 21188 19244 21244
rect 19244 21188 19248 21244
rect 19184 21184 19248 21188
rect 19264 21244 19328 21248
rect 19264 21188 19268 21244
rect 19268 21188 19324 21244
rect 19324 21188 19328 21244
rect 19264 21184 19328 21188
rect 3664 20700 3728 20704
rect 3664 20644 3668 20700
rect 3668 20644 3724 20700
rect 3724 20644 3728 20700
rect 3664 20640 3728 20644
rect 3744 20700 3808 20704
rect 3744 20644 3748 20700
rect 3748 20644 3804 20700
rect 3804 20644 3808 20700
rect 3744 20640 3808 20644
rect 3824 20700 3888 20704
rect 3824 20644 3828 20700
rect 3828 20644 3884 20700
rect 3884 20644 3888 20700
rect 3824 20640 3888 20644
rect 3904 20700 3968 20704
rect 3904 20644 3908 20700
rect 3908 20644 3964 20700
rect 3964 20644 3968 20700
rect 3904 20640 3968 20644
rect 19024 20156 19088 20160
rect 19024 20100 19028 20156
rect 19028 20100 19084 20156
rect 19084 20100 19088 20156
rect 19024 20096 19088 20100
rect 19104 20156 19168 20160
rect 19104 20100 19108 20156
rect 19108 20100 19164 20156
rect 19164 20100 19168 20156
rect 19104 20096 19168 20100
rect 19184 20156 19248 20160
rect 19184 20100 19188 20156
rect 19188 20100 19244 20156
rect 19244 20100 19248 20156
rect 19184 20096 19248 20100
rect 19264 20156 19328 20160
rect 19264 20100 19268 20156
rect 19268 20100 19324 20156
rect 19324 20100 19328 20156
rect 19264 20096 19328 20100
rect 3664 19612 3728 19616
rect 3664 19556 3668 19612
rect 3668 19556 3724 19612
rect 3724 19556 3728 19612
rect 3664 19552 3728 19556
rect 3744 19612 3808 19616
rect 3744 19556 3748 19612
rect 3748 19556 3804 19612
rect 3804 19556 3808 19612
rect 3744 19552 3808 19556
rect 3824 19612 3888 19616
rect 3824 19556 3828 19612
rect 3828 19556 3884 19612
rect 3884 19556 3888 19612
rect 3824 19552 3888 19556
rect 3904 19612 3968 19616
rect 3904 19556 3908 19612
rect 3908 19556 3964 19612
rect 3964 19556 3968 19612
rect 3904 19552 3968 19556
rect 19024 19068 19088 19072
rect 19024 19012 19028 19068
rect 19028 19012 19084 19068
rect 19084 19012 19088 19068
rect 19024 19008 19088 19012
rect 19104 19068 19168 19072
rect 19104 19012 19108 19068
rect 19108 19012 19164 19068
rect 19164 19012 19168 19068
rect 19104 19008 19168 19012
rect 19184 19068 19248 19072
rect 19184 19012 19188 19068
rect 19188 19012 19244 19068
rect 19244 19012 19248 19068
rect 19184 19008 19248 19012
rect 19264 19068 19328 19072
rect 19264 19012 19268 19068
rect 19268 19012 19324 19068
rect 19324 19012 19328 19068
rect 19264 19008 19328 19012
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 19024 17980 19088 17984
rect 19024 17924 19028 17980
rect 19028 17924 19084 17980
rect 19084 17924 19088 17980
rect 19024 17920 19088 17924
rect 19104 17980 19168 17984
rect 19104 17924 19108 17980
rect 19108 17924 19164 17980
rect 19164 17924 19168 17980
rect 19104 17920 19168 17924
rect 19184 17980 19248 17984
rect 19184 17924 19188 17980
rect 19188 17924 19244 17980
rect 19244 17924 19248 17980
rect 19184 17920 19248 17924
rect 19264 17980 19328 17984
rect 19264 17924 19268 17980
rect 19268 17924 19324 17980
rect 19324 17924 19328 17980
rect 19264 17920 19328 17924
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 19024 16892 19088 16896
rect 19024 16836 19028 16892
rect 19028 16836 19084 16892
rect 19084 16836 19088 16892
rect 19024 16832 19088 16836
rect 19104 16892 19168 16896
rect 19104 16836 19108 16892
rect 19108 16836 19164 16892
rect 19164 16836 19168 16892
rect 19104 16832 19168 16836
rect 19184 16892 19248 16896
rect 19184 16836 19188 16892
rect 19188 16836 19244 16892
rect 19244 16836 19248 16892
rect 19184 16832 19248 16836
rect 19264 16892 19328 16896
rect 19264 16836 19268 16892
rect 19268 16836 19324 16892
rect 19324 16836 19328 16892
rect 19264 16832 19328 16836
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 19024 15804 19088 15808
rect 19024 15748 19028 15804
rect 19028 15748 19084 15804
rect 19084 15748 19088 15804
rect 19024 15744 19088 15748
rect 19104 15804 19168 15808
rect 19104 15748 19108 15804
rect 19108 15748 19164 15804
rect 19164 15748 19168 15804
rect 19104 15744 19168 15748
rect 19184 15804 19248 15808
rect 19184 15748 19188 15804
rect 19188 15748 19244 15804
rect 19244 15748 19248 15804
rect 19184 15744 19248 15748
rect 19264 15804 19328 15808
rect 19264 15748 19268 15804
rect 19268 15748 19324 15804
rect 19324 15748 19328 15804
rect 19264 15744 19328 15748
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 19024 14716 19088 14720
rect 19024 14660 19028 14716
rect 19028 14660 19084 14716
rect 19084 14660 19088 14716
rect 19024 14656 19088 14660
rect 19104 14716 19168 14720
rect 19104 14660 19108 14716
rect 19108 14660 19164 14716
rect 19164 14660 19168 14716
rect 19104 14656 19168 14660
rect 19184 14716 19248 14720
rect 19184 14660 19188 14716
rect 19188 14660 19244 14716
rect 19244 14660 19248 14716
rect 19184 14656 19248 14660
rect 19264 14716 19328 14720
rect 19264 14660 19268 14716
rect 19268 14660 19324 14716
rect 19324 14660 19328 14716
rect 19264 14656 19328 14660
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 19024 13628 19088 13632
rect 19024 13572 19028 13628
rect 19028 13572 19084 13628
rect 19084 13572 19088 13628
rect 19024 13568 19088 13572
rect 19104 13628 19168 13632
rect 19104 13572 19108 13628
rect 19108 13572 19164 13628
rect 19164 13572 19168 13628
rect 19104 13568 19168 13572
rect 19184 13628 19248 13632
rect 19184 13572 19188 13628
rect 19188 13572 19244 13628
rect 19244 13572 19248 13628
rect 19184 13568 19248 13572
rect 19264 13628 19328 13632
rect 19264 13572 19268 13628
rect 19268 13572 19324 13628
rect 19324 13572 19328 13628
rect 19264 13568 19328 13572
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 19024 12540 19088 12544
rect 19024 12484 19028 12540
rect 19028 12484 19084 12540
rect 19084 12484 19088 12540
rect 19024 12480 19088 12484
rect 19104 12540 19168 12544
rect 19104 12484 19108 12540
rect 19108 12484 19164 12540
rect 19164 12484 19168 12540
rect 19104 12480 19168 12484
rect 19184 12540 19248 12544
rect 19184 12484 19188 12540
rect 19188 12484 19244 12540
rect 19244 12484 19248 12540
rect 19184 12480 19248 12484
rect 19264 12540 19328 12544
rect 19264 12484 19268 12540
rect 19268 12484 19324 12540
rect 19324 12484 19328 12540
rect 19264 12480 19328 12484
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 19024 11452 19088 11456
rect 19024 11396 19028 11452
rect 19028 11396 19084 11452
rect 19084 11396 19088 11452
rect 19024 11392 19088 11396
rect 19104 11452 19168 11456
rect 19104 11396 19108 11452
rect 19108 11396 19164 11452
rect 19164 11396 19168 11452
rect 19104 11392 19168 11396
rect 19184 11452 19248 11456
rect 19184 11396 19188 11452
rect 19188 11396 19244 11452
rect 19244 11396 19248 11452
rect 19184 11392 19248 11396
rect 19264 11452 19328 11456
rect 19264 11396 19268 11452
rect 19268 11396 19324 11452
rect 19324 11396 19328 11452
rect 19264 11392 19328 11396
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 19024 10364 19088 10368
rect 19024 10308 19028 10364
rect 19028 10308 19084 10364
rect 19084 10308 19088 10364
rect 19024 10304 19088 10308
rect 19104 10364 19168 10368
rect 19104 10308 19108 10364
rect 19108 10308 19164 10364
rect 19164 10308 19168 10364
rect 19104 10304 19168 10308
rect 19184 10364 19248 10368
rect 19184 10308 19188 10364
rect 19188 10308 19244 10364
rect 19244 10308 19248 10364
rect 19184 10304 19248 10308
rect 19264 10364 19328 10368
rect 19264 10308 19268 10364
rect 19268 10308 19324 10364
rect 19324 10308 19328 10364
rect 19264 10304 19328 10308
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 19024 9276 19088 9280
rect 19024 9220 19028 9276
rect 19028 9220 19084 9276
rect 19084 9220 19088 9276
rect 19024 9216 19088 9220
rect 19104 9276 19168 9280
rect 19104 9220 19108 9276
rect 19108 9220 19164 9276
rect 19164 9220 19168 9276
rect 19104 9216 19168 9220
rect 19184 9276 19248 9280
rect 19184 9220 19188 9276
rect 19188 9220 19244 9276
rect 19244 9220 19248 9276
rect 19184 9216 19248 9220
rect 19264 9276 19328 9280
rect 19264 9220 19268 9276
rect 19268 9220 19324 9276
rect 19324 9220 19328 9276
rect 19264 9216 19328 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 19024 8188 19088 8192
rect 19024 8132 19028 8188
rect 19028 8132 19084 8188
rect 19084 8132 19088 8188
rect 19024 8128 19088 8132
rect 19104 8188 19168 8192
rect 19104 8132 19108 8188
rect 19108 8132 19164 8188
rect 19164 8132 19168 8188
rect 19104 8128 19168 8132
rect 19184 8188 19248 8192
rect 19184 8132 19188 8188
rect 19188 8132 19244 8188
rect 19244 8132 19248 8188
rect 19184 8128 19248 8132
rect 19264 8188 19328 8192
rect 19264 8132 19268 8188
rect 19268 8132 19324 8188
rect 19324 8132 19328 8188
rect 19264 8128 19328 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 19024 7100 19088 7104
rect 19024 7044 19028 7100
rect 19028 7044 19084 7100
rect 19084 7044 19088 7100
rect 19024 7040 19088 7044
rect 19104 7100 19168 7104
rect 19104 7044 19108 7100
rect 19108 7044 19164 7100
rect 19164 7044 19168 7100
rect 19104 7040 19168 7044
rect 19184 7100 19248 7104
rect 19184 7044 19188 7100
rect 19188 7044 19244 7100
rect 19244 7044 19248 7100
rect 19184 7040 19248 7044
rect 19264 7100 19328 7104
rect 19264 7044 19268 7100
rect 19268 7044 19324 7100
rect 19324 7044 19328 7100
rect 19264 7040 19328 7044
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 19024 6012 19088 6016
rect 19024 5956 19028 6012
rect 19028 5956 19084 6012
rect 19084 5956 19088 6012
rect 19024 5952 19088 5956
rect 19104 6012 19168 6016
rect 19104 5956 19108 6012
rect 19108 5956 19164 6012
rect 19164 5956 19168 6012
rect 19104 5952 19168 5956
rect 19184 6012 19248 6016
rect 19184 5956 19188 6012
rect 19188 5956 19244 6012
rect 19244 5956 19248 6012
rect 19184 5952 19248 5956
rect 19264 6012 19328 6016
rect 19264 5956 19268 6012
rect 19268 5956 19324 6012
rect 19324 5956 19328 6012
rect 19264 5952 19328 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 19024 4924 19088 4928
rect 19024 4868 19028 4924
rect 19028 4868 19084 4924
rect 19084 4868 19088 4924
rect 19024 4864 19088 4868
rect 19104 4924 19168 4928
rect 19104 4868 19108 4924
rect 19108 4868 19164 4924
rect 19164 4868 19168 4924
rect 19104 4864 19168 4868
rect 19184 4924 19248 4928
rect 19184 4868 19188 4924
rect 19188 4868 19244 4924
rect 19244 4868 19248 4924
rect 19184 4864 19248 4868
rect 19264 4924 19328 4928
rect 19264 4868 19268 4924
rect 19268 4868 19324 4924
rect 19324 4868 19328 4924
rect 19264 4864 19328 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 19024 3836 19088 3840
rect 19024 3780 19028 3836
rect 19028 3780 19084 3836
rect 19084 3780 19088 3836
rect 19024 3776 19088 3780
rect 19104 3836 19168 3840
rect 19104 3780 19108 3836
rect 19108 3780 19164 3836
rect 19164 3780 19168 3836
rect 19104 3776 19168 3780
rect 19184 3836 19248 3840
rect 19184 3780 19188 3836
rect 19188 3780 19244 3836
rect 19244 3780 19248 3836
rect 19184 3776 19248 3780
rect 19264 3836 19328 3840
rect 19264 3780 19268 3836
rect 19268 3780 19324 3836
rect 19324 3780 19328 3836
rect 19264 3776 19328 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 19024 2748 19088 2752
rect 19024 2692 19028 2748
rect 19028 2692 19084 2748
rect 19084 2692 19088 2748
rect 19024 2688 19088 2692
rect 19104 2748 19168 2752
rect 19104 2692 19108 2748
rect 19108 2692 19164 2748
rect 19164 2692 19168 2748
rect 19104 2688 19168 2692
rect 19184 2748 19248 2752
rect 19184 2692 19188 2748
rect 19188 2692 19244 2748
rect 19244 2692 19248 2748
rect 19184 2688 19248 2692
rect 19264 2748 19328 2752
rect 19264 2692 19268 2748
rect 19268 2692 19324 2748
rect 19324 2692 19328 2748
rect 19264 2688 19328 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 19024 1660 19088 1664
rect 19024 1604 19028 1660
rect 19028 1604 19084 1660
rect 19084 1604 19088 1660
rect 19024 1600 19088 1604
rect 19104 1660 19168 1664
rect 19104 1604 19108 1660
rect 19108 1604 19164 1660
rect 19164 1604 19168 1660
rect 19104 1600 19168 1604
rect 19184 1660 19248 1664
rect 19184 1604 19188 1660
rect 19188 1604 19244 1660
rect 19244 1604 19248 1660
rect 19184 1600 19248 1604
rect 19264 1660 19328 1664
rect 19264 1604 19268 1660
rect 19268 1604 19324 1660
rect 19324 1604 19328 1660
rect 19264 1600 19328 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 19024 572 19088 576
rect 19024 516 19028 572
rect 19028 516 19084 572
rect 19084 516 19088 572
rect 19024 512 19088 516
rect 19104 572 19168 576
rect 19104 516 19108 572
rect 19108 516 19164 572
rect 19164 516 19168 572
rect 19104 512 19168 516
rect 19184 572 19248 576
rect 19184 516 19188 572
rect 19188 516 19244 572
rect 19244 516 19248 572
rect 19184 512 19248 516
rect 19264 572 19328 576
rect 19264 516 19268 572
rect 19268 516 19324 572
rect 19324 516 19328 572
rect 19264 512 19328 516
<< metal4 >>
rect 3700 23892 3940 23900
rect 3696 23440 3940 23892
rect 19050 23440 19260 23630
rect 3656 22880 3976 23440
rect 3656 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3976 22880
rect 3656 21792 3976 22816
rect 3656 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3976 21792
rect 3656 20704 3976 21728
rect 3656 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3976 20704
rect 3656 19616 3976 20640
rect 3656 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3976 19616
rect 3656 18528 3976 19552
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 3656 17440 3976 18464
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3656 15264 3976 16288
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3656 14176 3976 15200
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3656 12000 3976 13024
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 19016 23424 19336 23440
rect 19016 23360 19024 23424
rect 19088 23360 19104 23424
rect 19168 23360 19184 23424
rect 19248 23360 19264 23424
rect 19328 23360 19336 23424
rect 19016 22336 19336 23360
rect 19016 22272 19024 22336
rect 19088 22272 19104 22336
rect 19168 22272 19184 22336
rect 19248 22272 19264 22336
rect 19328 22272 19336 22336
rect 19016 21248 19336 22272
rect 19016 21184 19024 21248
rect 19088 21184 19104 21248
rect 19168 21184 19184 21248
rect 19248 21184 19264 21248
rect 19328 21184 19336 21248
rect 19016 20160 19336 21184
rect 19016 20096 19024 20160
rect 19088 20096 19104 20160
rect 19168 20096 19184 20160
rect 19248 20096 19264 20160
rect 19328 20096 19336 20160
rect 19016 19072 19336 20096
rect 19016 19008 19024 19072
rect 19088 19008 19104 19072
rect 19168 19008 19184 19072
rect 19248 19008 19264 19072
rect 19328 19008 19336 19072
rect 19016 17984 19336 19008
rect 19016 17920 19024 17984
rect 19088 17920 19104 17984
rect 19168 17920 19184 17984
rect 19248 17920 19264 17984
rect 19328 17920 19336 17984
rect 19016 16896 19336 17920
rect 19016 16832 19024 16896
rect 19088 16832 19104 16896
rect 19168 16832 19184 16896
rect 19248 16832 19264 16896
rect 19328 16832 19336 16896
rect 19016 15808 19336 16832
rect 19016 15744 19024 15808
rect 19088 15744 19104 15808
rect 19168 15744 19184 15808
rect 19248 15744 19264 15808
rect 19328 15744 19336 15808
rect 19016 14720 19336 15744
rect 19016 14656 19024 14720
rect 19088 14656 19104 14720
rect 19168 14656 19184 14720
rect 19248 14656 19264 14720
rect 19328 14656 19336 14720
rect 19016 13632 19336 14656
rect 19016 13568 19024 13632
rect 19088 13568 19104 13632
rect 19168 13568 19184 13632
rect 19248 13568 19264 13632
rect 19328 13568 19336 13632
rect 19016 12544 19336 13568
rect 19016 12480 19024 12544
rect 19088 12480 19104 12544
rect 19168 12480 19184 12544
rect 19248 12480 19264 12544
rect 19328 12480 19336 12544
rect 19016 11456 19336 12480
rect 19016 11392 19024 11456
rect 19088 11392 19104 11456
rect 19168 11392 19184 11456
rect 19248 11392 19264 11456
rect 19328 11392 19336 11456
rect 19016 10368 19336 11392
rect 19016 10304 19024 10368
rect 19088 10304 19104 10368
rect 19168 10304 19184 10368
rect 19248 10304 19264 10368
rect 19328 10304 19336 10368
rect 19016 9280 19336 10304
rect 19016 9216 19024 9280
rect 19088 9216 19104 9280
rect 19168 9216 19184 9280
rect 19248 9216 19264 9280
rect 19328 9216 19336 9280
rect 19016 8192 19336 9216
rect 19016 8128 19024 8192
rect 19088 8128 19104 8192
rect 19168 8128 19184 8192
rect 19248 8128 19264 8192
rect 19328 8128 19336 8192
rect 19016 7104 19336 8128
rect 19016 7040 19024 7104
rect 19088 7040 19104 7104
rect 19168 7040 19184 7104
rect 19248 7040 19264 7104
rect 19328 7040 19336 7104
rect 19016 6016 19336 7040
rect 19016 5952 19024 6016
rect 19088 5952 19104 6016
rect 19168 5952 19184 6016
rect 19248 5952 19264 6016
rect 19328 5952 19336 6016
rect 19016 4928 19336 5952
rect 19016 4864 19024 4928
rect 19088 4864 19104 4928
rect 19168 4864 19184 4928
rect 19248 4864 19264 4928
rect 19328 4864 19336 4928
rect 19016 3840 19336 4864
rect 19016 3776 19024 3840
rect 19088 3776 19104 3840
rect 19168 3776 19184 3840
rect 19248 3776 19264 3840
rect 19328 3776 19336 3840
rect 19016 2752 19336 3776
rect 19016 2688 19024 2752
rect 19088 2688 19104 2752
rect 19168 2688 19184 2752
rect 19248 2688 19264 2752
rect 19328 2688 19336 2752
rect 19016 1664 19336 2688
rect 19016 1600 19024 1664
rect 19088 1600 19104 1664
rect 19168 1600 19184 1664
rect 19248 1600 19264 1664
rect 19328 1600 19336 1664
rect 19016 576 19336 1600
rect 19016 512 19024 576
rect 19088 512 19104 576
rect 19168 512 19184 576
rect 19248 512 19264 576
rect 19328 512 19336 576
rect 19016 496 19336 512
rect 19020 320 19320 496
use sky130_fd_sc_hd__or4_2  _0501_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5980 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0502_
timestamp 1694700623
transform 1 0 8556 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0503_
timestamp 1694700623
transform 1 0 11684 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0504_
timestamp 1694700623
transform 1 0 15088 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0505_
timestamp 1694700623
transform 1 0 17296 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0506_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 19136 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0507_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 20424 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0508_
timestamp 1694700623
transform 1 0 21896 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0509_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 22540 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0510_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 21896 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0511_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 22080 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0512_
timestamp 1694700623
transform 1 0 5796 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0513_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4232 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0514_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3864 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0515_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 19412 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0516_
timestamp 1694700623
transform 1 0 18860 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0517_
timestamp 1694700623
transform 1 0 4692 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1694700623
transform -1 0 3956 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0519_
timestamp 1694700623
transform 1 0 4140 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0520_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4416 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0521_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4876 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0522_
timestamp 1694700623
transform 1 0 4784 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0523_
timestamp 1694700623
transform -1 0 4508 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0524_
timestamp 1694700623
transform 1 0 4968 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0525_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5796 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0526_
timestamp 1694700623
transform -1 0 6256 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0527_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5152 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0528_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5796 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0529_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4508 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0530_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5796 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _0531_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6440 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _0532_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 15548 0 1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__and3_1  _0533_
timestamp 1694700623
transform 1 0 7360 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0534_
timestamp 1694700623
transform -1 0 7360 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0535_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7084 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0536_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6532 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0537_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6532 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0538_
timestamp 1694700623
transform 1 0 6532 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0539_
timestamp 1694700623
transform -1 0 6716 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0540_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 14628 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0541_
timestamp 1694700623
transform -1 0 7728 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0542_
timestamp 1694700623
transform -1 0 6992 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0543_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _0544_
timestamp 1694700623
transform -1 0 10396 0 1 21216
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0545_
timestamp 1694700623
transform -1 0 5704 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0546_
timestamp 1694700623
transform -1 0 5612 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0547_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6532 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _0548_
timestamp 1694700623
transform 1 0 7452 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0549_
timestamp 1694700623
transform -1 0 7912 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0550_
timestamp 1694700623
transform -1 0 8740 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0551_
timestamp 1694700623
transform -1 0 7268 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0552_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6992 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0553_
timestamp 1694700623
transform 1 0 6992 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0554_
timestamp 1694700623
transform -1 0 6624 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0555_
timestamp 1694700623
transform 1 0 9016 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0556_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7912 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0557_
timestamp 1694700623
transform 1 0 7452 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0558_
timestamp 1694700623
transform 1 0 7820 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _0559_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 14168 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _0560_
timestamp 1694700623
transform 1 0 13524 0 -1 21216
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _0561_
timestamp 1694700623
transform -1 0 5796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _0562_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5796 0 -1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0563_
timestamp 1694700623
transform 1 0 4968 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0564_
timestamp 1694700623
transform -1 0 9844 0 -1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_2  _0565_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5612 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0566_
timestamp 1694700623
transform 1 0 6256 0 1 19040
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_1  _0567_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 9016 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0568_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7544 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0569_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 9016 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0570_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 8464 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0571_
timestamp 1694700623
transform 1 0 7360 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0572_
timestamp 1694700623
transform -1 0 8924 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0573_
timestamp 1694700623
transform -1 0 8648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0574_
timestamp 1694700623
transform -1 0 8832 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _0575_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7912 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0576_
timestamp 1694700623
transform -1 0 13984 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0577_
timestamp 1694700623
transform -1 0 16836 0 1 19040
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0578_
timestamp 1694700623
transform -1 0 5060 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0579_
timestamp 1694700623
transform 1 0 4600 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0580_
timestamp 1694700623
transform 1 0 5888 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_2  _0581_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4876 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0582_
timestamp 1694700623
transform 1 0 7452 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0583_
timestamp 1694700623
transform 1 0 8648 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0584_
timestamp 1694700623
transform 1 0 6992 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0585_
timestamp 1694700623
transform -1 0 9568 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0586_
timestamp 1694700623
transform 1 0 9292 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0587_
timestamp 1694700623
transform -1 0 10396 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0588_
timestamp 1694700623
transform -1 0 7176 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0589_
timestamp 1694700623
transform 1 0 9384 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0590_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 10120 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0591_
timestamp 1694700623
transform -1 0 10856 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0592_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9844 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0593_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 13064 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0594_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 13800 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_4  _0595_
timestamp 1694700623
transform 1 0 14812 0 1 21216
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_2  _0596_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4692 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__a2bb2o_1  _0597_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6532 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _0598_
timestamp 1694700623
transform 1 0 5796 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0599_
timestamp 1694700623
transform 1 0 9016 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_4  _0600_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 20424 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0601_
timestamp 1694700623
transform -1 0 17204 0 1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_1  _0602_
timestamp 1694700623
transform 1 0 6992 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0603_
timestamp 1694700623
transform 1 0 7728 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0604_
timestamp 1694700623
transform 1 0 9384 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0605_
timestamp 1694700623
transform 1 0 10672 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0606_
timestamp 1694700623
transform 1 0 9752 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0607_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9936 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0608_
timestamp 1694700623
transform -1 0 11500 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0609_
timestamp 1694700623
transform -1 0 11592 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0610_
timestamp 1694700623
transform 1 0 11040 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0611_
timestamp 1694700623
transform -1 0 10856 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0612_
timestamp 1694700623
transform 1 0 11132 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0613_
timestamp 1694700623
transform -1 0 11592 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0614_
timestamp 1694700623
transform 1 0 10580 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _0615_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10948 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _0616_
timestamp 1694700623
transform -1 0 20516 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0617_
timestamp 1694700623
transform 1 0 18124 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0618_
timestamp 1694700623
transform 1 0 18676 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0619_
timestamp 1694700623
transform -1 0 19872 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__o211a_1  _0620_
timestamp 1694700623
transform -1 0 6532 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _0621_
timestamp 1694700623
transform 1 0 13984 0 -1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _0622_
timestamp 1694700623
transform 1 0 6808 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0623_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6992 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0624_
timestamp 1694700623
transform -1 0 7544 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _0625_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6808 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0626_
timestamp 1694700623
transform 1 0 9016 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0627_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9844 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0628_
timestamp 1694700623
transform 1 0 10304 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0629_
timestamp 1694700623
transform 1 0 6532 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0630_
timestamp 1694700623
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0631_
timestamp 1694700623
transform 1 0 10948 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0632_
timestamp 1694700623
transform 1 0 11132 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0633_
timestamp 1694700623
transform 1 0 11316 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0634_
timestamp 1694700623
transform 1 0 11500 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0635_
timestamp 1694700623
transform 1 0 11776 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0636_
timestamp 1694700623
transform 1 0 12420 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0637_
timestamp 1694700623
transform 1 0 11960 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_4  _0638_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 18584 0 -1 22304
box -38 -48 1418 592
use sky130_fd_sc_hd__a21oi_2  _0639_
timestamp 1694700623
transform 1 0 15364 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0640_
timestamp 1694700623
transform 1 0 14904 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0641_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 17204 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0642_
timestamp 1694700623
transform -1 0 18124 0 1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_1  _0643_
timestamp 1694700623
transform -1 0 7636 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0644_
timestamp 1694700623
transform -1 0 8280 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0645_
timestamp 1694700623
transform 1 0 7820 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0646_
timestamp 1694700623
transform 1 0 9476 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0647_
timestamp 1694700623
transform 1 0 10028 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0648_
timestamp 1694700623
transform 1 0 10212 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0649_
timestamp 1694700623
transform 1 0 11224 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0650_
timestamp 1694700623
transform 1 0 12236 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0651_
timestamp 1694700623
transform 1 0 11592 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0652_
timestamp 1694700623
transform 1 0 11776 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0653_
timestamp 1694700623
transform -1 0 14720 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_1  _0654_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 12604 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0655_
timestamp 1694700623
transform 1 0 11776 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0656_
timestamp 1694700623
transform 1 0 12236 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0657_
timestamp 1694700623
transform 1 0 13524 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0658_
timestamp 1694700623
transform -1 0 14352 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0659_
timestamp 1694700623
transform 1 0 15180 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0660_
timestamp 1694700623
transform 1 0 11040 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0661_
timestamp 1694700623
transform -1 0 12972 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_4  _0662_
timestamp 1694700623
transform 1 0 16100 0 -1 22304
box -38 -48 1418 592
use sky130_fd_sc_hd__and3_1  _0663_
timestamp 1694700623
transform 1 0 13064 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0664_
timestamp 1694700623
transform 1 0 13064 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0665_
timestamp 1694700623
transform -1 0 12972 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0666_
timestamp 1694700623
transform -1 0 7820 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0667_
timestamp 1694700623
transform 1 0 8188 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0668_
timestamp 1694700623
transform 1 0 9568 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0669_
timestamp 1694700623
transform 1 0 11040 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _0670_
timestamp 1694700623
transform -1 0 10304 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0671_
timestamp 1694700623
transform 1 0 11592 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0672_
timestamp 1694700623
transform -1 0 13984 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0673_
timestamp 1694700623
transform -1 0 13984 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _0674_
timestamp 1694700623
transform 1 0 13156 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0675_
timestamp 1694700623
transform -1 0 14076 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0676_
timestamp 1694700623
transform 1 0 14168 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0677_
timestamp 1694700623
transform 1 0 14352 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1694700623
transform -1 0 13708 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0679_
timestamp 1694700623
transform -1 0 8188 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0680_
timestamp 1694700623
transform 1 0 7820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0681_
timestamp 1694700623
transform 1 0 8372 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _0682_
timestamp 1694700623
transform 1 0 9568 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0683_
timestamp 1694700623
transform 1 0 10396 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0684_
timestamp 1694700623
transform -1 0 11500 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0685_
timestamp 1694700623
transform 1 0 11316 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0686_
timestamp 1694700623
transform 1 0 13524 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0687_
timestamp 1694700623
transform 1 0 12420 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0688_
timestamp 1694700623
transform -1 0 14812 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0689_
timestamp 1694700623
transform 1 0 13800 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0690_
timestamp 1694700623
transform -1 0 10856 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_1  _0691_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 13064 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0692_
timestamp 1694700623
transform -1 0 12788 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0693_
timestamp 1694700623
transform -1 0 14720 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_1  _0694_
timestamp 1694700623
transform -1 0 13248 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0695_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 14076 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0696_
timestamp 1694700623
transform 1 0 14628 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0697_
timestamp 1694700623
transform 1 0 15180 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0698_
timestamp 1694700623
transform 1 0 15180 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0699_
timestamp 1694700623
transform -1 0 12972 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0700_
timestamp 1694700623
transform -1 0 12788 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0701_
timestamp 1694700623
transform 1 0 9660 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _0702_
timestamp 1694700623
transform 1 0 8188 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0703_
timestamp 1694700623
transform 1 0 10948 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0704_
timestamp 1694700623
transform 1 0 12236 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0705_
timestamp 1694700623
transform 1 0 14076 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0706_
timestamp 1694700623
transform -1 0 15272 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0707_
timestamp 1694700623
transform 1 0 14444 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0708_
timestamp 1694700623
transform 1 0 14904 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0709_
timestamp 1694700623
transform -1 0 16468 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0710_
timestamp 1694700623
transform -1 0 16284 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0711_
timestamp 1694700623
transform -1 0 4416 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0712_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5980 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0713_
timestamp 1694700623
transform 1 0 8280 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0714_
timestamp 1694700623
transform 1 0 10120 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0715_
timestamp 1694700623
transform 1 0 13340 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _0716_
timestamp 1694700623
transform -1 0 10948 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0717_
timestamp 1694700623
transform 1 0 14536 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0718_
timestamp 1694700623
transform -1 0 16744 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0719_
timestamp 1694700623
transform -1 0 12420 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0720_
timestamp 1694700623
transform -1 0 12236 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0721_
timestamp 1694700623
transform 1 0 15916 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0722_
timestamp 1694700623
transform -1 0 14168 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0723_
timestamp 1694700623
transform 1 0 13340 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0724_
timestamp 1694700623
transform -1 0 14260 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0725_
timestamp 1694700623
transform -1 0 16100 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0726_
timestamp 1694700623
transform 1 0 17296 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0727_
timestamp 1694700623
transform 1 0 16376 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0728_
timestamp 1694700623
transform -1 0 18216 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0729_
timestamp 1694700623
transform 1 0 16652 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0730_
timestamp 1694700623
transform 1 0 16100 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _0731_
timestamp 1694700623
transform -1 0 8188 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0732_
timestamp 1694700623
transform -1 0 18400 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0733_
timestamp 1694700623
transform 1 0 16100 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0734_
timestamp 1694700623
transform 1 0 10948 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0735_
timestamp 1694700623
transform -1 0 11868 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0736_
timestamp 1694700623
transform -1 0 18032 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0737_
timestamp 1694700623
transform -1 0 17480 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _0738_
timestamp 1694700623
transform 1 0 14720 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_2  _0739_
timestamp 1694700623
transform 1 0 15456 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0740_
timestamp 1694700623
transform 1 0 16468 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0741_
timestamp 1694700623
transform 1 0 15640 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0742_
timestamp 1694700623
transform -1 0 16836 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0743_
timestamp 1694700623
transform 1 0 16836 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1694700623
transform 1 0 17204 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0745_
timestamp 1694700623
transform -1 0 16744 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0746_
timestamp 1694700623
transform -1 0 17572 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0747_
timestamp 1694700623
transform -1 0 16008 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0748_
timestamp 1694700623
transform -1 0 16100 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0749_
timestamp 1694700623
transform 1 0 16836 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0750_
timestamp 1694700623
transform -1 0 17756 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0751_
timestamp 1694700623
transform 1 0 17572 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0752_
timestamp 1694700623
transform 1 0 17756 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0753_
timestamp 1694700623
transform 1 0 17848 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0754_
timestamp 1694700623
transform 1 0 17480 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0755_
timestamp 1694700623
transform 1 0 18676 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0756_
timestamp 1694700623
transform 1 0 18032 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0757_
timestamp 1694700623
transform -1 0 19320 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0758_
timestamp 1694700623
transform -1 0 18584 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0759_
timestamp 1694700623
transform -1 0 17848 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0760_
timestamp 1694700623
transform 1 0 18308 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0761_
timestamp 1694700623
transform -1 0 17572 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0762_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14168 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0763_
timestamp 1694700623
transform -1 0 17940 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0764_
timestamp 1694700623
transform 1 0 17388 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0765_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 16652 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0766_
timestamp 1694700623
transform 1 0 18124 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0767_
timestamp 1694700623
transform 1 0 18676 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1694700623
transform 1 0 19596 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0769_
timestamp 1694700623
transform -1 0 18584 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0770_
timestamp 1694700623
transform -1 0 20148 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0771_
timestamp 1694700623
transform 1 0 20700 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1694700623
transform -1 0 20700 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0773_
timestamp 1694700623
transform -1 0 20240 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0774_
timestamp 1694700623
transform 1 0 19320 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0775_
timestamp 1694700623
transform -1 0 18584 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0776_
timestamp 1694700623
transform -1 0 20424 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0777_
timestamp 1694700623
transform -1 0 19320 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0778_
timestamp 1694700623
transform 1 0 18676 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0779_
timestamp 1694700623
transform 1 0 19044 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0780_
timestamp 1694700623
transform -1 0 19872 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1694700623
transform -1 0 18768 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0782_
timestamp 1694700623
transform 1 0 19504 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0783_
timestamp 1694700623
transform 1 0 19504 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0784_
timestamp 1694700623
transform 1 0 18676 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1694700623
transform -1 0 19596 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0786_
timestamp 1694700623
transform 1 0 20148 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0787_
timestamp 1694700623
transform -1 0 19504 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0788_
timestamp 1694700623
transform -1 0 19504 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1694700623
transform 1 0 19136 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0790_
timestamp 1694700623
transform -1 0 20148 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0791_
timestamp 1694700623
transform 1 0 20700 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0792_
timestamp 1694700623
transform 1 0 21344 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0793_
timestamp 1694700623
transform -1 0 22448 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0794_
timestamp 1694700623
transform -1 0 23000 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0795_
timestamp 1694700623
transform -1 0 22264 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0796_
timestamp 1694700623
transform 1 0 21528 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0797_
timestamp 1694700623
transform 1 0 22080 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0798_
timestamp 1694700623
transform -1 0 22632 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0799_
timestamp 1694700623
transform 1 0 20240 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0800_
timestamp 1694700623
transform -1 0 20884 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0801_
timestamp 1694700623
transform 1 0 20056 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0802_
timestamp 1694700623
transform 1 0 20332 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1694700623
transform -1 0 21988 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0804_
timestamp 1694700623
transform 1 0 20700 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0805_
timestamp 1694700623
transform 1 0 21160 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0806_
timestamp 1694700623
transform 1 0 21252 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0807_
timestamp 1694700623
transform -1 0 21988 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _0808_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 20608 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0809_
timestamp 1694700623
transform 1 0 21896 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0810_
timestamp 1694700623
transform -1 0 22264 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0811_
timestamp 1694700623
transform 1 0 22264 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0812_
timestamp 1694700623
transform -1 0 22540 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _0813_
timestamp 1694700623
transform 1 0 21712 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0814_
timestamp 1694700623
transform -1 0 21160 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0815_
timestamp 1694700623
transform 1 0 21160 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0816_
timestamp 1694700623
transform 1 0 20884 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0817_
timestamp 1694700623
transform -1 0 21344 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0818_
timestamp 1694700623
transform 1 0 21344 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0819_
timestamp 1694700623
transform 1 0 21252 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0820_
timestamp 1694700623
transform -1 0 23092 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0821_
timestamp 1694700623
transform -1 0 21160 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0822_
timestamp 1694700623
transform -1 0 21528 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0823_
timestamp 1694700623
transform -1 0 21712 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _0824_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6440 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0825_
timestamp 1694700623
transform 1 0 5796 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0826_
timestamp 1694700623
transform 1 0 5520 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0827_
timestamp 1694700623
transform -1 0 5520 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0828_
timestamp 1694700623
transform 1 0 5796 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0829_
timestamp 1694700623
transform -1 0 6624 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0830_
timestamp 1694700623
transform 1 0 5060 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp 1694700623
transform -1 0 6164 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0832_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6164 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0833_
timestamp 1694700623
transform 1 0 6624 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0834_
timestamp 1694700623
transform 1 0 7084 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0835_
timestamp 1694700623
transform -1 0 7820 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0836_
timestamp 1694700623
transform 1 0 7820 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0837_
timestamp 1694700623
transform -1 0 8188 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0838_
timestamp 1694700623
transform 1 0 7544 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0839_
timestamp 1694700623
transform 1 0 9844 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0840_
timestamp 1694700623
transform 1 0 8832 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0841_
timestamp 1694700623
transform -1 0 9016 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0842_
timestamp 1694700623
transform 1 0 8188 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0843_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9016 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0844_
timestamp 1694700623
transform 1 0 8004 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0845_
timestamp 1694700623
transform 1 0 9568 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0846_
timestamp 1694700623
transform 1 0 10028 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0847_
timestamp 1694700623
transform 1 0 10304 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0848_
timestamp 1694700623
transform -1 0 11684 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0849_
timestamp 1694700623
transform -1 0 11224 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0850_
timestamp 1694700623
transform 1 0 11408 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0851_
timestamp 1694700623
transform 1 0 10580 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0852_
timestamp 1694700623
transform 1 0 10764 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0853_
timestamp 1694700623
transform 1 0 12052 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0854_
timestamp 1694700623
transform 1 0 10948 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0855_
timestamp 1694700623
transform 1 0 12604 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0856_
timestamp 1694700623
transform 1 0 13524 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0857_
timestamp 1694700623
transform -1 0 14260 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0858_
timestamp 1694700623
transform 1 0 14260 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0859_
timestamp 1694700623
transform 1 0 14720 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0860_
timestamp 1694700623
transform -1 0 14812 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0861_
timestamp 1694700623
transform -1 0 14260 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0862_
timestamp 1694700623
transform 1 0 13616 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0863_
timestamp 1694700623
transform 1 0 14168 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0864_
timestamp 1694700623
transform 1 0 14720 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0865_
timestamp 1694700623
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0866_
timestamp 1694700623
transform 1 0 15824 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0867_
timestamp 1694700623
transform -1 0 16284 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0868_
timestamp 1694700623
transform -1 0 17388 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0869_
timestamp 1694700623
transform -1 0 16836 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0870_
timestamp 1694700623
transform 1 0 16468 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0871_
timestamp 1694700623
transform 1 0 16284 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0872_
timestamp 1694700623
transform 1 0 17112 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0873_
timestamp 1694700623
transform 1 0 17756 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0874_
timestamp 1694700623
transform 1 0 16928 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 1694700623
transform 1 0 18124 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0876_
timestamp 1694700623
transform 1 0 18676 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0877_
timestamp 1694700623
transform 1 0 18676 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0878_
timestamp 1694700623
transform 1 0 19320 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0879_
timestamp 1694700623
transform 1 0 19596 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0880_
timestamp 1694700623
transform 1 0 19964 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0881_
timestamp 1694700623
transform 1 0 18676 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0882_
timestamp 1694700623
transform 1 0 19964 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0883_
timestamp 1694700623
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0884_
timestamp 1694700623
transform -1 0 21712 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0885_
timestamp 1694700623
transform -1 0 21068 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0886_
timestamp 1694700623
transform 1 0 20884 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0887_
timestamp 1694700623
transform -1 0 21712 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0888_
timestamp 1694700623
transform 1 0 21252 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0889_
timestamp 1694700623
transform 1 0 20792 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0890_
timestamp 1694700623
transform 1 0 22356 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0891_
timestamp 1694700623
transform -1 0 22356 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0892_
timestamp 1694700623
transform 1 0 21252 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0893_
timestamp 1694700623
transform -1 0 23000 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0894_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 21528 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0895_
timestamp 1694700623
transform 1 0 19412 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0896_
timestamp 1694700623
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0897_
timestamp 1694700623
transform 1 0 20516 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0898_
timestamp 1694700623
transform 1 0 21344 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 1694700623
transform -1 0 22172 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0900_
timestamp 1694700623
transform -1 0 22356 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0901_
timestamp 1694700623
transform -1 0 22816 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0902_
timestamp 1694700623
transform 1 0 20700 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0903_
timestamp 1694700623
transform -1 0 6072 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0904_
timestamp 1694700623
transform -1 0 5060 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0905_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7728 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0906_
timestamp 1694700623
transform 1 0 5796 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0907_
timestamp 1694700623
transform 1 0 4600 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0908_
timestamp 1694700623
transform -1 0 20976 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 1694700623
transform -1 0 6992 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0910_
timestamp 1694700623
transform -1 0 7728 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 1694700623
transform -1 0 4600 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0912_
timestamp 1694700623
transform 1 0 5796 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0913_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5704 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0914_
timestamp 1694700623
transform -1 0 5060 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0915_
timestamp 1694700623
transform 1 0 5244 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0916_
timestamp 1694700623
transform 1 0 4876 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0917_
timestamp 1694700623
transform -1 0 7544 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0918_
timestamp 1694700623
transform 1 0 6532 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0919_
timestamp 1694700623
transform -1 0 5704 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0920_
timestamp 1694700623
transform -1 0 4324 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0921_
timestamp 1694700623
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0922_
timestamp 1694700623
transform 1 0 22724 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0923_
timestamp 1694700623
transform 1 0 5888 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0924_
timestamp 1694700623
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0925_
timestamp 1694700623
transform -1 0 7728 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0926_
timestamp 1694700623
transform -1 0 7360 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0927_
timestamp 1694700623
transform 1 0 7820 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0928_
timestamp 1694700623
transform -1 0 8280 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0929_
timestamp 1694700623
transform -1 0 8280 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0930_
timestamp 1694700623
transform -1 0 7636 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0931_
timestamp 1694700623
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0932_
timestamp 1694700623
transform 1 0 8372 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0933_
timestamp 1694700623
transform 1 0 8740 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0934_
timestamp 1694700623
transform -1 0 10580 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0935_
timestamp 1694700623
transform -1 0 9384 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0936_
timestamp 1694700623
transform -1 0 10304 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0937_
timestamp 1694700623
transform 1 0 10304 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0938_
timestamp 1694700623
transform 1 0 9384 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1694700623
transform -1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0940_
timestamp 1694700623
transform 1 0 10764 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0941_
timestamp 1694700623
transform -1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0942_
timestamp 1694700623
transform -1 0 11776 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0943_
timestamp 1694700623
transform -1 0 12972 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0944_
timestamp 1694700623
transform -1 0 12788 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0945_
timestamp 1694700623
transform 1 0 12972 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0946_
timestamp 1694700623
transform -1 0 15456 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0947_
timestamp 1694700623
transform -1 0 14904 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0948_
timestamp 1694700623
transform -1 0 12788 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0949_
timestamp 1694700623
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0950_
timestamp 1694700623
transform -1 0 14996 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0951_
timestamp 1694700623
transform -1 0 14260 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0952_
timestamp 1694700623
transform 1 0 17572 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0953_
timestamp 1694700623
transform -1 0 16008 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0954_
timestamp 1694700623
transform -1 0 17480 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0955_
timestamp 1694700623
transform -1 0 15640 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0956_
timestamp 1694700623
transform -1 0 16284 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0957_
timestamp 1694700623
transform -1 0 16376 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0958_
timestamp 1694700623
transform 1 0 16284 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0959_
timestamp 1694700623
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1694700623
transform 1 0 16376 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0961_
timestamp 1694700623
transform 1 0 20240 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0962_
timestamp 1694700623
transform -1 0 18124 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0963_
timestamp 1694700623
transform 1 0 18124 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0964_
timestamp 1694700623
transform -1 0 19964 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0965_
timestamp 1694700623
transform -1 0 20240 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1694700623
transform -1 0 18124 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0967_
timestamp 1694700623
transform 1 0 18768 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0968_
timestamp 1694700623
transform 1 0 19964 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0969_
timestamp 1694700623
transform -1 0 19964 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0970_
timestamp 1694700623
transform -1 0 21160 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0971_
timestamp 1694700623
transform -1 0 20976 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0972_
timestamp 1694700623
transform -1 0 22080 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0973_
timestamp 1694700623
transform 1 0 21068 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0974_
timestamp 1694700623
transform 1 0 20516 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0975_
timestamp 1694700623
transform -1 0 22356 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0976_
timestamp 1694700623
transform -1 0 21804 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0977_
timestamp 1694700623
transform -1 0 20700 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0978_
timestamp 1694700623
transform 1 0 22540 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0979_
timestamp 1694700623
transform -1 0 22172 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0980_
timestamp 1694700623
transform -1 0 20700 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0981_
timestamp 1694700623
transform -1 0 22448 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0982_
timestamp 1694700623
transform 1 0 21344 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0983_
timestamp 1694700623
transform 1 0 20700 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0984_
timestamp 1694700623
transform -1 0 22724 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0985_
timestamp 1694700623
transform -1 0 22632 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0986_
timestamp 1694700623
transform -1 0 22172 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0987_
timestamp 1694700623
transform -1 0 21712 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0988_
timestamp 1694700623
transform -1 0 19320 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0989_
timestamp 1694700623
transform 1 0 18768 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0990_
timestamp 1694700623
transform -1 0 18860 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1694700623
transform -1 0 18400 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1694700623
transform -1 0 19228 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0993_
timestamp 1694700623
transform 1 0 17572 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0994_
timestamp 1694700623
transform -1 0 18584 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0995_
timestamp 1694700623
transform -1 0 20700 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0996_
timestamp 1694700623
transform 1 0 20884 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0997_
timestamp 1694700623
transform 1 0 19872 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1694700623
transform 1 0 20240 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0999_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 19780 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1000_
timestamp 1694700623
transform 1 0 20148 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1001_
timestamp 1694700623
transform -1 0 22080 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1002_
timestamp 1694700623
transform -1 0 21436 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1003_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4232 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1694700623
transform 1 0 4324 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1694700623
transform 1 0 4508 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1694700623
transform 1 0 4232 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1694700623
transform 1 0 4876 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1694700623
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1694700623
transform -1 0 9844 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1694700623
transform 1 0 9384 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1694700623
transform -1 0 12420 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1694700623
transform 1 0 11500 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1694700623
transform -1 0 14996 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1694700623
transform 1 0 13708 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1694700623
transform 1 0 14536 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1694700623
transform 1 0 16100 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1694700623
transform 1 0 16284 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1694700623
transform 1 0 16744 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1694700623
transform 1 0 18676 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1694700623
transform -1 0 19872 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1694700623
transform 1 0 19688 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1694700623
transform -1 0 23092 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1694700623
transform 1 0 21160 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1694700623
transform 1 0 21252 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1694700623
transform 1 0 5796 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1694700623
transform -1 0 5704 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1694700623
transform 1 0 5060 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1694700623
transform 1 0 4968 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1694700623
transform 1 0 4232 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1694700623
transform 1 0 4324 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1694700623
transform -1 0 7268 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1694700623
transform 1 0 6348 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1694700623
transform 1 0 7452 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1694700623
transform -1 0 9292 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1694700623
transform 1 0 9384 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1694700623
transform -1 0 11500 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1694700623
transform -1 0 12420 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1694700623
transform 1 0 12512 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1694700623
transform 1 0 12788 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1694700623
transform 1 0 13524 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1694700623
transform 1 0 15548 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1694700623
transform 1 0 16100 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1694700623
transform 1 0 16100 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1694700623
transform 1 0 18676 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1694700623
transform 1 0 18124 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1694700623
transform -1 0 19688 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1694700623
transform 1 0 21252 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1694700623
transform -1 0 22448 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1694700623
transform -1 0 22540 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1694700623
transform 1 0 21252 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1694700623
transform -1 0 22908 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1694700623
transform 1 0 21436 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1694700623
transform 1 0 18676 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1694700623
transform 1 0 18032 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1694700623
transform 1 0 19964 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1694700623
transform 1 0 19688 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1694700623
transform 1 0 21252 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 9016 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  fanout13 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 17204 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1694700623
transform 1 0 5152 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout15
timestamp 1694700623
transform -1 0 11776 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout16
timestamp 1694700623
transform 1 0 20792 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout17
timestamp 1694700623
transform -1 0 9660 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp 1694700623
transform -1 0 14628 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 1694700623
transform 1 0 13156 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1694700623
transform -1 0 22540 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 1694700623
transform -1 0 23000 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 1694700623
transform 1 0 22724 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout23 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 22172 0 1 7072
box -38 -48 958 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1694700623
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1694700623
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1694700623
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1694700623
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1694700623
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1694700623
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1694700623
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1694700623
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1694700623
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1694700623
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1694700623
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1694700623
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1694700623
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1694700623
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1694700623
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1694700623
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1694700623
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1694700623
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1694700623
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1694700623
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1694700623
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1694700623
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_237 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 22356 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1694700623
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1694700623
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1694700623
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1694700623
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1694700623
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1694700623
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1694700623
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1694700623
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1694700623
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1694700623
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1694700623
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1694700623
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1694700623
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1694700623
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1694700623
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1694700623
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1694700623
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1694700623
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1694700623
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1694700623
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1694700623
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1694700623
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1694700623
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_237
timestamp 1694700623
transform 1 0 22356 0 -1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1694700623
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1694700623
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1694700623
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1694700623
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1694700623
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1694700623
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1694700623
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1694700623
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1694700623
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1694700623
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1694700623
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1694700623
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1694700623
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1694700623
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1694700623
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1694700623
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1694700623
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1694700623
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1694700623
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1694700623
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1694700623
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1694700623
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1694700623
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1694700623
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1694700623
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1694700623
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1694700623
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1694700623
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1694700623
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1694700623
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1694700623
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1694700623
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1694700623
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1694700623
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1694700623
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1694700623
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1694700623
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1694700623
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1694700623
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1694700623
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1694700623
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1694700623
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1694700623
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1694700623
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1694700623
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1694700623
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1694700623
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1694700623
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1694700623
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1694700623
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_237
timestamp 1694700623
transform 1 0 22356 0 -1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1694700623
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1694700623
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1694700623
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1694700623
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1694700623
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1694700623
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1694700623
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1694700623
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1694700623
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1694700623
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1694700623
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1694700623
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1694700623
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1694700623
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1694700623
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1694700623
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1694700623
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1694700623
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1694700623
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1694700623
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1694700623
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1694700623
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1694700623
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1694700623
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1694700623
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1694700623
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1694700623
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1694700623
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1694700623
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1694700623
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1694700623
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1694700623
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1694700623
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1694700623
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1694700623
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1694700623
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1694700623
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1694700623
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1694700623
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1694700623
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1694700623
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1694700623
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1694700623
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1694700623
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1694700623
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1694700623
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1694700623
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1694700623
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1694700623
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1694700623
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_237
timestamp 1694700623
transform 1 0 22356 0 -1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1694700623
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1694700623
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1694700623
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1694700623
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1694700623
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1694700623
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1694700623
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1694700623
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1694700623
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1694700623
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1694700623
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1694700623
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1694700623
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1694700623
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1694700623
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1694700623
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1694700623
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1694700623
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1694700623
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1694700623
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1694700623
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1694700623
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1694700623
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1694700623
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_233 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 21988 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1694700623
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1694700623
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1694700623
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1694700623
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1694700623
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1694700623
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_63
timestamp 1694700623
transform 1 0 6348 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_75
timestamp 1694700623
transform 1 0 7452 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_87
timestamp 1694700623
transform 1 0 8556 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_99
timestamp 1694700623
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1694700623
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1694700623
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1694700623
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1694700623
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1694700623
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1694700623
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1694700623
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1694700623
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1694700623
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1694700623
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_205
timestamp 1694700623
transform 1 0 19412 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_213
timestamp 1694700623
transform 1 0 20148 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1694700623
transform 1 0 20516 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1694700623
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1694700623
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_237
timestamp 1694700623
transform 1 0 22356 0 -1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1694700623
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1694700623
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1694700623
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1694700623
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_41
timestamp 1694700623
transform 1 0 4324 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_45
timestamp 1694700623
transform 1 0 4692 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1694700623
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1694700623
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1694700623
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1694700623
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1694700623
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1694700623
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1694700623
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1694700623
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1694700623
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1694700623
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1694700623
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1694700623
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1694700623
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1694700623
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1694700623
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_197
timestamp 1694700623
transform 1 0 18676 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_201
timestamp 1694700623
transform 1 0 19044 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_209
timestamp 1694700623
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_230
timestamp 1694700623
transform 1 0 21712 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_242
timestamp 1694700623
transform 1 0 22816 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1694700623
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1694700623
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1694700623
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_39
timestamp 1694700623
transform 1 0 4140 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_78
timestamp 1694700623
transform 1 0 7728 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_90
timestamp 1694700623
transform 1 0 8832 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_102
timestamp 1694700623
transform 1 0 9936 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1694700623
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1694700623
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1694700623
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1694700623
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1694700623
transform 1 0 14260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1694700623
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1694700623
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1694700623
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_181
timestamp 1694700623
transform 1 0 17204 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_189
timestamp 1694700623
transform 1 0 17940 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_206
timestamp 1694700623
transform 1 0 19504 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_225
timestamp 1694700623
transform 1 0 21252 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_243
timestamp 1694700623
transform 1 0 22908 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1694700623
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1694700623
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1694700623
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1694700623
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_78
timestamp 1694700623
transform 1 0 7728 0 1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1694700623
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1694700623
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1694700623
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1694700623
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1694700623
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1694700623
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1694700623
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1694700623
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1694700623
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_177
timestamp 1694700623
transform 1 0 16836 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_244
timestamp 1694700623
transform 1 0 23000 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1694700623
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1694700623
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1694700623
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_39
timestamp 1694700623
transform 1 0 4140 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_45
timestamp 1694700623
transform 1 0 4692 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_70
timestamp 1694700623
transform 1 0 6992 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_74
timestamp 1694700623
transform 1 0 7360 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_91
timestamp 1694700623
transform 1 0 8924 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_95
timestamp 1694700623
transform 1 0 9292 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_116
timestamp 1694700623
transform 1 0 11224 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_128
timestamp 1694700623
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1694700623
transform 1 0 14260 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1694700623
transform 1 0 15364 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1694700623
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_172
timestamp 1694700623
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_184
timestamp 1694700623
transform 1 0 17480 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_190
timestamp 1694700623
transform 1 0 18032 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_204
timestamp 1694700623
transform 1 0 19320 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1694700623
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_225
timestamp 1694700623
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_242
timestamp 1694700623
transform 1 0 22816 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1694700623
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1694700623
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1694700623
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1694700623
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1694700623
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_53
timestamp 1694700623
transform 1 0 5428 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_60
timestamp 1694700623
transform 1 0 6072 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_72
timestamp 1694700623
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_122
timestamp 1694700623
transform 1 0 11776 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_130
timestamp 1694700623
transform 1 0 12512 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_157
timestamp 1694700623
transform 1 0 14996 0 1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_179
timestamp 1694700623
transform 1 0 17020 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_191
timestamp 1694700623
transform 1 0 18124 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1694700623
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_197
timestamp 1694700623
transform 1 0 18676 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_203
timestamp 1694700623
transform 1 0 19228 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_219
timestamp 1694700623
transform 1 0 20700 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_225
timestamp 1694700623
transform 1 0 21252 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1694700623
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1694700623
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1694700623
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1694700623
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1694700623
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1694700623
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_57
timestamp 1694700623
transform 1 0 5796 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_99
timestamp 1694700623
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_162
timestamp 1694700623
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_189
timestamp 1694700623
transform 1 0 17940 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_201
timestamp 1694700623
transform 1 0 19044 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_213
timestamp 1694700623
transform 1 0 20148 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_221
timestamp 1694700623
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_225
timestamp 1694700623
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_243
timestamp 1694700623
transform 1 0 22908 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1694700623
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1694700623
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1694700623
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1694700623
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_41
timestamp 1694700623
transform 1 0 4324 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_55
timestamp 1694700623
transform 1 0 5612 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_65
timestamp 1694700623
transform 1 0 6532 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_69
timestamp 1694700623
transform 1 0 6900 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_93
timestamp 1694700623
transform 1 0 9108 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_109
timestamp 1694700623
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_123
timestamp 1694700623
transform 1 0 11868 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_129
timestamp 1694700623
transform 1 0 12420 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1694700623
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1694700623
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1694700623
transform 1 0 14996 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_188
timestamp 1694700623
transform 1 0 17848 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_213
timestamp 1694700623
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_241
timestamp 1694700623
transform 1 0 22724 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1694700623
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1694700623
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1694700623
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_39
timestamp 1694700623
transform 1 0 4140 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_73
timestamp 1694700623
transform 1 0 7268 0 -1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_84
timestamp 1694700623
transform 1 0 8280 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_96
timestamp 1694700623
transform 1 0 9384 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_108
timestamp 1694700623
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1694700623
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1694700623
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_141
timestamp 1694700623
transform 1 0 13524 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1694700623
transform 1 0 14260 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1694700623
transform 1 0 15364 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1694700623
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_185
timestamp 1694700623
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 1694700623
transform 1 0 20976 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1694700623
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1694700623
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1694700623
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_29
timestamp 1694700623
transform 1 0 3220 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_37
timestamp 1694700623
transform 1 0 3956 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_76
timestamp 1694700623
transform 1 0 7544 0 1 9248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1694700623
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1694700623
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_109
timestamp 1694700623
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_131
timestamp 1694700623
transform 1 0 12604 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1694700623
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_155
timestamp 1694700623
transform 1 0 14812 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_167
timestamp 1694700623
transform 1 0 15916 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_171
timestamp 1694700623
transform 1 0 16284 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_175
timestamp 1694700623
transform 1 0 16652 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_187
timestamp 1694700623
transform 1 0 17756 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_197
timestamp 1694700623
transform 1 0 18676 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_242
timestamp 1694700623
transform 1 0 22816 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1694700623
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1694700623
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1694700623
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_39
timestamp 1694700623
transform 1 0 4140 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_47
timestamp 1694700623
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_65
timestamp 1694700623
transform 1 0 6532 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_77
timestamp 1694700623
transform 1 0 7636 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_97
timestamp 1694700623
transform 1 0 9476 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_110
timestamp 1694700623
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_116
timestamp 1694700623
transform 1 0 11224 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_128
timestamp 1694700623
transform 1 0 12328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_140
timestamp 1694700623
transform 1 0 13432 0 -1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_154
timestamp 1694700623
transform 1 0 14720 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1694700623
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1694700623
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 1694700623
transform 1 0 17204 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_189
timestamp 1694700623
transform 1 0 17940 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_211
timestamp 1694700623
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_219
timestamp 1694700623
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_225
timestamp 1694700623
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_235
timestamp 1694700623
transform 1 0 22172 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_243
timestamp 1694700623
transform 1 0 22908 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1694700623
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1694700623
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1694700623
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1694700623
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_41
timestamp 1694700623
transform 1 0 4324 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_49
timestamp 1694700623
transform 1 0 5060 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_69
timestamp 1694700623
transform 1 0 6900 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_104
timestamp 1694700623
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_128
timestamp 1694700623
transform 1 0 12328 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_134
timestamp 1694700623
transform 1 0 12880 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1694700623
transform 1 0 13524 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_157
timestamp 1694700623
transform 1 0 14996 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_165
timestamp 1694700623
transform 1 0 15732 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_193
timestamp 1694700623
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1694700623
transform 1 0 18676 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_209
timestamp 1694700623
transform 1 0 19780 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_217
timestamp 1694700623
transform 1 0 20516 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_222
timestamp 1694700623
transform 1 0 20976 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_237
timestamp 1694700623
transform 1 0 22356 0 1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1694700623
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1694700623
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1694700623
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_39
timestamp 1694700623
transform 1 0 4140 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_47
timestamp 1694700623
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_69
timestamp 1694700623
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_94
timestamp 1694700623
transform 1 0 9200 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_106
timestamp 1694700623
transform 1 0 10304 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_135
timestamp 1694700623
transform 1 0 12972 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_143
timestamp 1694700623
transform 1 0 13708 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_149
timestamp 1694700623
transform 1 0 14260 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_153
timestamp 1694700623
transform 1 0 14628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_160
timestamp 1694700623
transform 1 0 15272 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_172
timestamp 1694700623
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_177
timestamp 1694700623
transform 1 0 16836 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_189
timestamp 1694700623
transform 1 0 17940 0 -1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_204
timestamp 1694700623
transform 1 0 19320 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_216
timestamp 1694700623
transform 1 0 20424 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_241
timestamp 1694700623
transform 1 0 22724 0 -1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1694700623
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1694700623
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1694700623
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1694700623
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_41
timestamp 1694700623
transform 1 0 4324 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_49
timestamp 1694700623
transform 1 0 5060 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_66
timestamp 1694700623
transform 1 0 6624 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_78
timestamp 1694700623
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1694700623
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1694700623
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1694700623
transform 1 0 9476 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_109
timestamp 1694700623
transform 1 0 10580 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_120
timestamp 1694700623
transform 1 0 11592 0 1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_127
timestamp 1694700623
transform 1 0 12236 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1694700623
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_157
timestamp 1694700623
transform 1 0 14996 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_165
timestamp 1694700623
transform 1 0 15732 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_183
timestamp 1694700623
transform 1 0 17388 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1694700623
transform 1 0 18492 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_217
timestamp 1694700623
transform 1 0 20516 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_221
timestamp 1694700623
transform 1 0 20884 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_238
timestamp 1694700623
transform 1 0 22448 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_244
timestamp 1694700623
transform 1 0 23000 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1694700623
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1694700623
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1694700623
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_39
timestamp 1694700623
transform 1 0 4140 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_45
timestamp 1694700623
transform 1 0 4692 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1694700623
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1694700623
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_69
timestamp 1694700623
transform 1 0 6900 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_81
timestamp 1694700623
transform 1 0 8004 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_90
timestamp 1694700623
transform 1 0 8832 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_138
timestamp 1694700623
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_162
timestamp 1694700623
transform 1 0 15456 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_169
timestamp 1694700623
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_177
timestamp 1694700623
transform 1 0 16836 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_184
timestamp 1694700623
transform 1 0 17480 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_190
timestamp 1694700623
transform 1 0 18032 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_194
timestamp 1694700623
transform 1 0 18400 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_206
timestamp 1694700623
transform 1 0 19504 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_218
timestamp 1694700623
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1694700623
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1694700623
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1694700623
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_29
timestamp 1694700623
transform 1 0 3220 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_37
timestamp 1694700623
transform 1 0 3956 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_59
timestamp 1694700623
transform 1 0 5980 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_67
timestamp 1694700623
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_101
timestamp 1694700623
transform 1 0 9844 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_112
timestamp 1694700623
transform 1 0 10856 0 1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_122
timestamp 1694700623
transform 1 0 11776 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_134
timestamp 1694700623
transform 1 0 12880 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_162
timestamp 1694700623
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_173
timestamp 1694700623
transform 1 0 16468 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_181
timestamp 1694700623
transform 1 0 17204 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1694700623
transform 1 0 17940 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1694700623
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_204
timestamp 1694700623
transform 1 0 19320 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_216
timestamp 1694700623
transform 1 0 20424 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_244
timestamp 1694700623
transform 1 0 23000 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1694700623
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1694700623
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_27
timestamp 1694700623
transform 1 0 3036 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_33
timestamp 1694700623
transform 1 0 3588 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_66
timestamp 1694700623
transform 1 0 6624 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_78
timestamp 1694700623
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_91
timestamp 1694700623
transform 1 0 8924 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_99
timestamp 1694700623
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_108
timestamp 1694700623
transform 1 0 10488 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_120
timestamp 1694700623
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_129
timestamp 1694700623
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_141
timestamp 1694700623
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_149
timestamp 1694700623
transform 1 0 14260 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_185
timestamp 1694700623
transform 1 0 17572 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_197
timestamp 1694700623
transform 1 0 18676 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_201
timestamp 1694700623
transform 1 0 19044 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_214
timestamp 1694700623
transform 1 0 20240 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_220
timestamp 1694700623
transform 1 0 20792 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_230
timestamp 1694700623
transform 1 0 21712 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_242
timestamp 1694700623
transform 1 0 22816 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1694700623
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1694700623
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1694700623
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1694700623
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_57
timestamp 1694700623
transform 1 0 5796 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_69
timestamp 1694700623
transform 1 0 6900 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_73
timestamp 1694700623
transform 1 0 7268 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1694700623
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_88
timestamp 1694700623
transform 1 0 8648 0 1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_101
timestamp 1694700623
transform 1 0 9844 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_113
timestamp 1694700623
transform 1 0 10948 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_123
timestamp 1694700623
transform 1 0 11868 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_135
timestamp 1694700623
transform 1 0 12972 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1694700623
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_155
timestamp 1694700623
transform 1 0 14812 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_171
timestamp 1694700623
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_192
timestamp 1694700623
transform 1 0 18216 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_197
timestamp 1694700623
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_208
timestamp 1694700623
transform 1 0 19688 0 1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_228
timestamp 1694700623
transform 1 0 21528 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_240
timestamp 1694700623
transform 1 0 22632 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_244
timestamp 1694700623
transform 1 0 23000 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1694700623
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1694700623
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1694700623
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_39
timestamp 1694700623
transform 1 0 4140 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1694700623
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_57
timestamp 1694700623
transform 1 0 5796 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_86
timestamp 1694700623
transform 1 0 8464 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_94
timestamp 1694700623
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_120
timestamp 1694700623
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_136
timestamp 1694700623
transform 1 0 13064 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_147
timestamp 1694700623
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_159
timestamp 1694700623
transform 1 0 15180 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1694700623
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1694700623
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_190
timestamp 1694700623
transform 1 0 18032 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_210
timestamp 1694700623
transform 1 0 19872 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_218
timestamp 1694700623
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_240
timestamp 1694700623
transform 1 0 22632 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_244
timestamp 1694700623
transform 1 0 23000 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1694700623
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1694700623
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1694700623
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1694700623
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_41
timestamp 1694700623
transform 1 0 4324 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_63
timestamp 1694700623
transform 1 0 6348 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_95
timestamp 1694700623
transform 1 0 9292 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_107
timestamp 1694700623
transform 1 0 10396 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_115
timestamp 1694700623
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_131
timestamp 1694700623
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1694700623
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_154
timestamp 1694700623
transform 1 0 14720 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_166
timestamp 1694700623
transform 1 0 15824 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_170
timestamp 1694700623
transform 1 0 16192 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_192
timestamp 1694700623
transform 1 0 18216 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_216
timestamp 1694700623
transform 1 0 20424 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_239
timestamp 1694700623
transform 1 0 22540 0 1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1694700623
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1694700623
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1694700623
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_39
timestamp 1694700623
transform 1 0 4140 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_78
timestamp 1694700623
transform 1 0 7728 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_89
timestamp 1694700623
transform 1 0 8740 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_97
timestamp 1694700623
transform 1 0 9476 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_107
timestamp 1694700623
transform 1 0 10396 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1694700623
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_119
timestamp 1694700623
transform 1 0 11500 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_131
timestamp 1694700623
transform 1 0 12604 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_147
timestamp 1694700623
transform 1 0 14076 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_160
timestamp 1694700623
transform 1 0 15272 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_169
timestamp 1694700623
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_187
timestamp 1694700623
transform 1 0 17756 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_195
timestamp 1694700623
transform 1 0 18492 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_216
timestamp 1694700623
transform 1 0 20424 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_241
timestamp 1694700623
transform 1 0 22724 0 -1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1694700623
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1694700623
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1694700623
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1694700623
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_41
timestamp 1694700623
transform 1 0 4324 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_45
timestamp 1694700623
transform 1 0 4692 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_71
timestamp 1694700623
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_80
timestamp 1694700623
transform 1 0 7912 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_85
timestamp 1694700623
transform 1 0 8372 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_93
timestamp 1694700623
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_108
timestamp 1694700623
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_123
timestamp 1694700623
transform 1 0 11868 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_135
timestamp 1694700623
transform 1 0 12972 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1694700623
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_141
timestamp 1694700623
transform 1 0 13524 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_169
timestamp 1694700623
transform 1 0 16100 0 1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_184
timestamp 1694700623
transform 1 0 17480 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1694700623
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1694700623
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_221
timestamp 1694700623
transform 1 0 20884 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_229
timestamp 1694700623
transform 1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1694700623
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1694700623
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1694700623
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1694700623
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1694700623
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1694700623
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_57
timestamp 1694700623
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_68
timestamp 1694700623
transform 1 0 6808 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_80
timestamp 1694700623
transform 1 0 7912 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_92
timestamp 1694700623
transform 1 0 9016 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_106
timestamp 1694700623
transform 1 0 10304 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_122
timestamp 1694700623
transform 1 0 11776 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_160
timestamp 1694700623
transform 1 0 15272 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_169
timestamp 1694700623
transform 1 0 16100 0 -1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_185
timestamp 1694700623
transform 1 0 17572 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_204
timestamp 1694700623
transform 1 0 19320 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_216
timestamp 1694700623
transform 1 0 20424 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_241
timestamp 1694700623
transform 1 0 22724 0 -1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1694700623
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1694700623
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1694700623
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1694700623
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1694700623
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1694700623
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1694700623
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1694700623
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1694700623
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_85
timestamp 1694700623
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_95
timestamp 1694700623
transform 1 0 9292 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_112
timestamp 1694700623
transform 1 0 10856 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_129
timestamp 1694700623
transform 1 0 12420 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_137
timestamp 1694700623
transform 1 0 13156 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_141
timestamp 1694700623
transform 1 0 13524 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_155
timestamp 1694700623
transform 1 0 14812 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_163
timestamp 1694700623
transform 1 0 15548 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_174
timestamp 1694700623
transform 1 0 16560 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_189
timestamp 1694700623
transform 1 0 17940 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_204
timestamp 1694700623
transform 1 0 19320 0 1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1694700623
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1694700623
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1694700623
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_39
timestamp 1694700623
transform 1 0 4140 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_43
timestamp 1694700623
transform 1 0 4508 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1694700623
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1694700623
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_70
timestamp 1694700623
transform 1 0 6992 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1694700623
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1694700623
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1694700623
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_137
timestamp 1694700623
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_154
timestamp 1694700623
transform 1 0 14720 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1694700623
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_176
timestamp 1694700623
transform 1 0 16744 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_188
timestamp 1694700623
transform 1 0 17848 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_194
timestamp 1694700623
transform 1 0 18400 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_210
timestamp 1694700623
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_228
timestamp 1694700623
transform 1 0 21528 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1694700623
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1694700623
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1694700623
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_29
timestamp 1694700623
transform 1 0 3220 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_35
timestamp 1694700623
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_43
timestamp 1694700623
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_68
timestamp 1694700623
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_82
timestamp 1694700623
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_92
timestamp 1694700623
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_104
timestamp 1694700623
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_113
timestamp 1694700623
transform 1 0 10948 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_149
timestamp 1694700623
transform 1 0 14260 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_153
timestamp 1694700623
transform 1 0 14628 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_160
timestamp 1694700623
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_184
timestamp 1694700623
transform 1 0 17480 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1694700623
transform 1 0 18676 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_209
timestamp 1694700623
transform 1 0 19780 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_239
timestamp 1694700623
transform 1 0 22540 0 1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1694700623
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1694700623
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1694700623
transform 1 0 3036 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1694700623
transform 1 0 4140 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1694700623
transform 1 0 5244 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1694700623
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_78
timestamp 1694700623
transform 1 0 7728 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_82
timestamp 1694700623
transform 1 0 8096 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_90
timestamp 1694700623
transform 1 0 8832 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_98
timestamp 1694700623
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_129
timestamp 1694700623
transform 1 0 12420 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_137
timestamp 1694700623
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1694700623
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1694700623
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_181
timestamp 1694700623
transform 1 0 17204 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_188
timestamp 1694700623
transform 1 0 17848 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_192
timestamp 1694700623
transform 1 0 18216 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_209
timestamp 1694700623
transform 1 0 19780 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_215
timestamp 1694700623
transform 1 0 20332 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1694700623
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_229
timestamp 1694700623
transform 1 0 21620 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_233
timestamp 1694700623
transform 1 0 21988 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_240
timestamp 1694700623
transform 1 0 22632 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_244
timestamp 1694700623
transform 1 0 23000 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1694700623
transform 1 0 828 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1694700623
transform 1 0 1932 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1694700623
transform 1 0 3036 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1694700623
transform 1 0 3220 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_41
timestamp 1694700623
transform 1 0 4324 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_45
timestamp 1694700623
transform 1 0 4692 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_93
timestamp 1694700623
transform 1 0 9108 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_101
timestamp 1694700623
transform 1 0 9844 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_123
timestamp 1694700623
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1694700623
transform 1 0 12788 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1694700623
transform 1 0 13340 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_154
timestamp 1694700623
transform 1 0 14720 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_213
timestamp 1694700623
transform 1 0 20148 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_240
timestamp 1694700623
transform 1 0 22632 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_244
timestamp 1694700623
transform 1 0 23000 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1694700623
transform 1 0 828 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1694700623
transform 1 0 1932 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1694700623
transform 1 0 3036 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_39
timestamp 1694700623
transform 1 0 4140 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_79
timestamp 1694700623
transform 1 0 7820 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_83
timestamp 1694700623
transform 1 0 8188 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_97
timestamp 1694700623
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1694700623
transform 1 0 10764 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_116
timestamp 1694700623
transform 1 0 11224 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_135
timestamp 1694700623
transform 1 0 12972 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_150
timestamp 1694700623
transform 1 0 14352 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_162
timestamp 1694700623
transform 1 0 15456 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_182
timestamp 1694700623
transform 1 0 17296 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_188
timestamp 1694700623
transform 1 0 17848 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_195
timestamp 1694700623
transform 1 0 18492 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1694700623
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_217
timestamp 1694700623
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_225
timestamp 1694700623
transform 1 0 21252 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_229
timestamp 1694700623
transform 1 0 21620 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_233
timestamp 1694700623
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1694700623
transform 1 0 828 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1694700623
transform 1 0 1932 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1694700623
transform 1 0 3036 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_29
timestamp 1694700623
transform 1 0 3220 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_37
timestamp 1694700623
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_47
timestamp 1694700623
transform 1 0 4876 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_57
timestamp 1694700623
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_65
timestamp 1694700623
transform 1 0 6532 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_69
timestamp 1694700623
transform 1 0 6900 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_76
timestamp 1694700623
transform 1 0 7544 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1694700623
transform 1 0 8188 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1694700623
transform 1 0 8372 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1694700623
transform 1 0 9476 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1694700623
transform 1 0 10580 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_121
timestamp 1694700623
transform 1 0 11684 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_129
timestamp 1694700623
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_135
timestamp 1694700623
transform 1 0 12972 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1694700623
transform 1 0 13340 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_146
timestamp 1694700623
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_194
timestamp 1694700623
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_202
timestamp 1694700623
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_214
timestamp 1694700623
transform 1 0 20240 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_220
timestamp 1694700623
transform 1 0 20792 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_240
timestamp 1694700623
transform 1 0 22632 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_244
timestamp 1694700623
transform 1 0 23000 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1694700623
transform 1 0 828 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1694700623
transform 1 0 1932 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1694700623
transform 1 0 3036 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_46
timestamp 1694700623
transform 1 0 4784 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_52
timestamp 1694700623
transform 1 0 5336 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_65
timestamp 1694700623
transform 1 0 6532 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_96
timestamp 1694700623
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1694700623
transform 1 0 10764 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_119
timestamp 1694700623
transform 1 0 11500 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_127
timestamp 1694700623
transform 1 0 12236 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_135
timestamp 1694700623
transform 1 0 12972 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_163
timestamp 1694700623
transform 1 0 15548 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1694700623
transform 1 0 15916 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_185
timestamp 1694700623
transform 1 0 17572 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_197
timestamp 1694700623
transform 1 0 18676 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_201
timestamp 1694700623
transform 1 0 19044 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1694700623
transform 1 0 19412 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_217
timestamp 1694700623
transform 1 0 20516 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_233
timestamp 1694700623
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1694700623
transform 1 0 828 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1694700623
transform 1 0 1932 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1694700623
transform 1 0 3036 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1694700623
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1694700623
transform 1 0 4324 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1694700623
transform 1 0 5428 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_65
timestamp 1694700623
transform 1 0 6532 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_74
timestamp 1694700623
transform 1 0 7360 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_113
timestamp 1694700623
transform 1 0 10948 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_181
timestamp 1694700623
transform 1 0 17204 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1694700623
transform 1 0 18308 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_213
timestamp 1694700623
transform 1 0 20148 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_240
timestamp 1694700623
transform 1 0 22632 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_244
timestamp 1694700623
transform 1 0 23000 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1694700623
transform 1 0 828 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1694700623
transform 1 0 1932 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1694700623
transform 1 0 3036 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_39
timestamp 1694700623
transform 1 0 4140 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_47
timestamp 1694700623
transform 1 0 4876 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_61
timestamp 1694700623
transform 1 0 6164 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1694700623
transform 1 0 10764 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_113
timestamp 1694700623
transform 1 0 10948 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_221
timestamp 1694700623
transform 1 0 20884 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_244
timestamp 1694700623
transform 1 0 23000 0 -1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1694700623
transform 1 0 828 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1694700623
transform 1 0 1932 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1694700623
transform 1 0 3036 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1694700623
transform 1 0 3220 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_41
timestamp 1694700623
transform 1 0 4324 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_53
timestamp 1694700623
transform 1 0 5428 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_64
timestamp 1694700623
transform 1 0 6440 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1694700623
transform 1 0 8188 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_85
timestamp 1694700623
transform 1 0 8372 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_89
timestamp 1694700623
transform 1 0 8740 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_135
timestamp 1694700623
transform 1 0 12972 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1694700623
transform 1 0 13340 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_217
timestamp 1694700623
transform 1 0 20516 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_236
timestamp 1694700623
transform 1 0 22264 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_244
timestamp 1694700623
transform 1 0 23000 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_3
timestamp 1694700623
transform 1 0 828 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_11
timestamp 1694700623
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_16
timestamp 1694700623
transform 1 0 2024 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_29
timestamp 1694700623
transform 1 0 3220 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_41
timestamp 1694700623
transform 1 0 4324 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1694700623
transform 1 0 5244 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1694700623
transform 1 0 5612 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_61
timestamp 1694700623
transform 1 0 6164 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_69
timestamp 1694700623
transform 1 0 6900 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_74
timestamp 1694700623
transform 1 0 7360 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_83
timestamp 1694700623
transform 1 0 8188 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_85
timestamp 1694700623
transform 1 0 8372 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_97
timestamp 1694700623
transform 1 0 9476 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1694700623
transform 1 0 10764 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_124
timestamp 1694700623
transform 1 0 11960 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_136
timestamp 1694700623
transform 1 0 13064 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_147
timestamp 1694700623
transform 1 0 14076 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_155
timestamp 1694700623
transform 1 0 14812 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_189
timestamp 1694700623
transform 1 0 17940 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_195
timestamp 1694700623
transform 1 0 18492 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_200
timestamp 1694700623
transform 1 0 18952 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_204
timestamp 1694700623
transform 1 0 19320 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_222
timestamp 1694700623
transform 1 0 20976 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1694700623
transform 1 0 21252 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_243
timestamp 1694700623
transform 1 0 22908 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1694700623
transform -1 0 23092 0 1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input2 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 23092 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1694700623
transform 1 0 1748 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1694700623
transform 1 0 4692 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1694700623
transform 1 0 7636 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input6 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10948 0 -1 23392
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input7
timestamp 1694700623
transform 1 0 13524 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1694700623
transform 1 0 17664 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1694700623
transform 1 0 19412 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1694700623
transform 1 0 22356 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap12
timestamp 1694700623
transform 1 0 14628 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_42
timestamp 1694700623
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 23368 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_43
timestamp 1694700623
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 23368 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_44
timestamp 1694700623
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_45
timestamp 1694700623
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 23368 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_46
timestamp 1694700623
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 23368 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_47
timestamp 1694700623
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 23368 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_48
timestamp 1694700623
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 23368 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_49
timestamp 1694700623
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 23368 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_50
timestamp 1694700623
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 23368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_51
timestamp 1694700623
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 23368 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_52
timestamp 1694700623
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 23368 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_53
timestamp 1694700623
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 23368 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_54
timestamp 1694700623
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 23368 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_55
timestamp 1694700623
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 23368 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_56
timestamp 1694700623
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 23368 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_57
timestamp 1694700623
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1694700623
transform -1 0 23368 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_58
timestamp 1694700623
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1694700623
transform -1 0 23368 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_59
timestamp 1694700623
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1694700623
transform -1 0 23368 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_60
timestamp 1694700623
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1694700623
transform -1 0 23368 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_61
timestamp 1694700623
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1694700623
transform -1 0 23368 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_62
timestamp 1694700623
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1694700623
transform -1 0 23368 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_63
timestamp 1694700623
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1694700623
transform -1 0 23368 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_64
timestamp 1694700623
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1694700623
transform -1 0 23368 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_65
timestamp 1694700623
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1694700623
transform -1 0 23368 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_66
timestamp 1694700623
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1694700623
transform -1 0 23368 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_67
timestamp 1694700623
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1694700623
transform -1 0 23368 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_68
timestamp 1694700623
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1694700623
transform -1 0 23368 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_69
timestamp 1694700623
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1694700623
transform -1 0 23368 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_70
timestamp 1694700623
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1694700623
transform -1 0 23368 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_71
timestamp 1694700623
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1694700623
transform -1 0 23368 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_72
timestamp 1694700623
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1694700623
transform -1 0 23368 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_73
timestamp 1694700623
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1694700623
transform -1 0 23368 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_74
timestamp 1694700623
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1694700623
transform -1 0 23368 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_75
timestamp 1694700623
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1694700623
transform -1 0 23368 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_76
timestamp 1694700623
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1694700623
transform -1 0 23368 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_77
timestamp 1694700623
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1694700623
transform -1 0 23368 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_78
timestamp 1694700623
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1694700623
transform -1 0 23368 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_79
timestamp 1694700623
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1694700623
transform -1 0 23368 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_80
timestamp 1694700623
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1694700623
transform -1 0 23368 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_81
timestamp 1694700623
transform 1 0 552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1694700623
transform -1 0 23368 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_82
timestamp 1694700623
transform 1 0 552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1694700623
transform -1 0 23368 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_83
timestamp 1694700623
transform 1 0 552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1694700623
transform -1 0 23368 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1694700623
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1694700623
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1694700623
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1694700623
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_89
timestamp 1694700623
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_90
timestamp 1694700623
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_91
timestamp 1694700623
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1694700623
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1694700623
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_94
timestamp 1694700623
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_95
timestamp 1694700623
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1694700623
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1694700623
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1694700623
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1694700623
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1694700623
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1694700623
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1694700623
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1694700623
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_104
timestamp 1694700623
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1694700623
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1694700623
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1694700623
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_108
timestamp 1694700623
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_109
timestamp 1694700623
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_110
timestamp 1694700623
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1694700623
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_112
timestamp 1694700623
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_113
timestamp 1694700623
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_114
timestamp 1694700623
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_115
timestamp 1694700623
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1694700623
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_117
timestamp 1694700623
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_118
timestamp 1694700623
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_119
timestamp 1694700623
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1694700623
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1694700623
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1694700623
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_123
timestamp 1694700623
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1694700623
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1694700623
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1694700623
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1694700623
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1694700623
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1694700623
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1694700623
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1694700623
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp 1694700623
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp 1694700623
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1694700623
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1694700623
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_136
timestamp 1694700623
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_137
timestamp 1694700623
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_138
timestamp 1694700623
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1694700623
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_140
timestamp 1694700623
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_141
timestamp 1694700623
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_142
timestamp 1694700623
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_143
timestamp 1694700623
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_144
timestamp 1694700623
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_145
timestamp 1694700623
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_146
timestamp 1694700623
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_147
timestamp 1694700623
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_148
timestamp 1694700623
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_149
timestamp 1694700623
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_150
timestamp 1694700623
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_151
timestamp 1694700623
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_152
timestamp 1694700623
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_153
timestamp 1694700623
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_154
timestamp 1694700623
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_155
timestamp 1694700623
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp 1694700623
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_157
timestamp 1694700623
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_158
timestamp 1694700623
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_159
timestamp 1694700623
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp 1694700623
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp 1694700623
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_162
timestamp 1694700623
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_163
timestamp 1694700623
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp 1694700623
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp 1694700623
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_166
timestamp 1694700623
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_167
timestamp 1694700623
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp 1694700623
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp 1694700623
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_170
timestamp 1694700623
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_171
timestamp 1694700623
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp 1694700623
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp 1694700623
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_174
timestamp 1694700623
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_175
timestamp 1694700623
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_176
timestamp 1694700623
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp 1694700623
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_178
timestamp 1694700623
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_179
timestamp 1694700623
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_180
timestamp 1694700623
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_181
timestamp 1694700623
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_182
timestamp 1694700623
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_183
timestamp 1694700623
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_184
timestamp 1694700623
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_185
timestamp 1694700623
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_186
timestamp 1694700623
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_187
timestamp 1694700623
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_188
timestamp 1694700623
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_189
timestamp 1694700623
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_190
timestamp 1694700623
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_191
timestamp 1694700623
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_192
timestamp 1694700623
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_193
timestamp 1694700623
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_194
timestamp 1694700623
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_195
timestamp 1694700623
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_196
timestamp 1694700623
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_197
timestamp 1694700623
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_198
timestamp 1694700623
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_199
timestamp 1694700623
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_200
timestamp 1694700623
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_201
timestamp 1694700623
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_202
timestamp 1694700623
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_203
timestamp 1694700623
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_204
timestamp 1694700623
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_205
timestamp 1694700623
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_206
timestamp 1694700623
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_207
timestamp 1694700623
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_208
timestamp 1694700623
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_209
timestamp 1694700623
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_210
timestamp 1694700623
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_211
timestamp 1694700623
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_212
timestamp 1694700623
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_213
timestamp 1694700623
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_214
timestamp 1694700623
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_215
timestamp 1694700623
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_216
timestamp 1694700623
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_217
timestamp 1694700623
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_218
timestamp 1694700623
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_219
timestamp 1694700623
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_220
timestamp 1694700623
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_221
timestamp 1694700623
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_222
timestamp 1694700623
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_223
timestamp 1694700623
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_224
timestamp 1694700623
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_225
timestamp 1694700623
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_226
timestamp 1694700623
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_227
timestamp 1694700623
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_228
timestamp 1694700623
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_229
timestamp 1694700623
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_230
timestamp 1694700623
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_231
timestamp 1694700623
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_232
timestamp 1694700623
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_233
timestamp 1694700623
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_234
timestamp 1694700623
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_235
timestamp 1694700623
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_236
timestamp 1694700623
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_237
timestamp 1694700623
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_238
timestamp 1694700623
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_239
timestamp 1694700623
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_240
timestamp 1694700623
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_241
timestamp 1694700623
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_242
timestamp 1694700623
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_243
timestamp 1694700623
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_244
timestamp 1694700623
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_245
timestamp 1694700623
transform 1 0 10856 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_246
timestamp 1694700623
transform 1 0 16008 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_247
timestamp 1694700623
transform 1 0 21160 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_248
timestamp 1694700623
transform 1 0 3128 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_249
timestamp 1694700623
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_250
timestamp 1694700623
transform 1 0 13432 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_251
timestamp 1694700623
transform 1 0 18584 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_252
timestamp 1694700623
transform 1 0 3128 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_253
timestamp 1694700623
transform 1 0 5704 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_254
timestamp 1694700623
transform 1 0 8280 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_255
timestamp 1694700623
transform 1 0 10856 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_256
timestamp 1694700623
transform 1 0 13432 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_257
timestamp 1694700623
transform 1 0 16008 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_258
timestamp 1694700623
transform 1 0 18584 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_259
timestamp 1694700623
transform 1 0 21160 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire11
timestamp 1694700623
transform -1 0 13432 0 -1 15776
box -38 -48 314 592
<< labels >>
flabel metal4 s 19016 496 19336 23440 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3656 496 3976 23440 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 23600 3816 24000 3936 0 FreeSans 480 0 0 0 clk_in
port 2 nsew signal input
flabel metal3 s 23600 19592 24000 19712 0 FreeSans 480 0 0 0 clk_out
port 3 nsew signal tristate
flabel metal3 s 23600 11704 24000 11824 0 FreeSans 480 0 0 0 nrst
port 4 nsew signal input
flabel metal2 s 1674 23600 1730 24000 0 FreeSans 224 90 0 0 scale[0]
port 5 nsew signal input
flabel metal2 s 4618 23600 4674 24000 0 FreeSans 224 90 0 0 scale[1]
port 6 nsew signal input
flabel metal2 s 7562 23600 7618 24000 0 FreeSans 224 90 0 0 scale[2]
port 7 nsew signal input
flabel metal2 s 10506 23600 10562 24000 0 FreeSans 224 90 0 0 scale[3]
port 8 nsew signal input
flabel metal2 s 13450 23600 13506 24000 0 FreeSans 224 90 0 0 scale[4]
port 9 nsew signal input
flabel metal2 s 16394 23600 16450 24000 0 FreeSans 224 90 0 0 scale[5]
port 10 nsew signal input
flabel metal2 s 19338 23600 19394 24000 0 FreeSans 224 90 0 0 scale[6]
port 11 nsew signal input
flabel metal2 s 22282 23600 22338 24000 0 FreeSans 224 90 0 0 scale[7]
port 12 nsew signal input
rlabel metal1 11960 23392 11960 23392 0 VGND
rlabel metal1 11960 22848 11960 22848 0 VPWR
rlabel metal1 4354 13430 4354 13430 0 _0000_
rlabel metal1 4002 13498 4002 13498 0 _0001_
rlabel metal1 4630 12682 4630 12682 0 _0002_
rlabel metal1 4871 15606 4871 15606 0 _0003_
rlabel metal1 5423 14926 5423 14926 0 _0004_
rlabel metal1 7309 12682 7309 12682 0 _0005_
rlabel metal1 8928 12750 8928 12750 0 _0006_
rlabel metal1 9793 12342 9793 12342 0 _0007_
rlabel metal1 11826 12342 11826 12342 0 _0008_
rlabel metal1 11909 11254 11909 11254 0 _0009_
rlabel metal1 14776 11662 14776 11662 0 _0010_
rlabel metal1 13830 12342 13830 12342 0 _0011_
rlabel metal1 15180 12954 15180 12954 0 _0012_
rlabel metal1 16314 13430 16314 13430 0 _0013_
rlabel via1 16601 14926 16601 14926 0 _0014_
rlabel metal1 16964 13838 16964 13838 0 _0015_
rlabel metal1 18752 14858 18752 14858 0 _0016_
rlabel metal1 19887 14518 19887 14518 0 _0017_
rlabel metal1 20189 17102 20189 17102 0 _0018_
rlabel metal1 22544 17782 22544 17782 0 _0019_
rlabel metal1 21380 17102 21380 17102 0 _0020_
rlabel metal1 21615 16694 21615 16694 0 _0021_
rlabel metal1 5382 5338 5382 5338 0 _0022_
rlabel metal1 5704 4794 5704 4794 0 _0023_
rlabel metal1 4952 5066 4952 5066 0 _0024_
rlabel via1 5280 6222 5280 6222 0 _0025_
rlabel metal1 4733 9010 4733 9010 0 _0026_
rlabel metal1 4446 9418 4446 9418 0 _0027_
rlabel metal1 6348 8602 6348 8602 0 _0028_
rlabel metal1 6987 7990 6987 7990 0 _0029_
rlabel metal1 7666 6902 7666 6902 0 _0030_
rlabel metal1 8878 7514 8878 7514 0 _0031_
rlabel metal2 9706 7174 9706 7174 0 _0032_
rlabel metal2 11178 7106 11178 7106 0 _0033_
rlabel metal2 11730 7718 11730 7718 0 _0034_
rlabel viali 12829 6902 12829 6902 0 _0035_
rlabel metal1 12910 7990 12910 7990 0 _0036_
rlabel metal2 14122 7106 14122 7106 0 _0037_
rlabel via1 15865 7310 15865 7310 0 _0038_
rlabel metal1 16376 6970 16376 6970 0 _0039_
rlabel metal1 16463 9078 16463 9078 0 _0040_
rlabel metal1 18896 8398 18896 8398 0 _0041_
rlabel metal1 18338 9078 18338 9078 0 _0042_
rlabel metal1 19611 10166 19611 10166 0 _0043_
rlabel metal1 21242 11186 21242 11186 0 _0044_
rlabel metal2 22310 11186 22310 11186 0 _0045_
rlabel metal1 22463 9418 22463 9418 0 _0046_
rlabel metal1 21334 9010 21334 9010 0 _0047_
rlabel viali 22590 7922 22590 7922 0 _0048_
rlabel metal1 21712 5338 21712 5338 0 _0049_
rlabel metal1 18896 6222 18896 6222 0 _0050_
rlabel metal1 18441 5814 18441 5814 0 _0051_
rlabel metal2 20286 4930 20286 4930 0 _0052_
rlabel metal1 20097 5814 20097 5814 0 _0053_
rlabel metal2 21390 15334 21390 15334 0 _0054_
rlabel metal1 7268 10982 7268 10982 0 _0055_
rlabel metal1 9752 10574 9752 10574 0 _0056_
rlabel metal1 12834 10608 12834 10608 0 _0057_
rlabel metal2 17250 12478 17250 12478 0 _0058_
rlabel metal1 18814 12852 18814 12852 0 _0059_
rlabel metal1 20194 13430 20194 13430 0 _0060_
rlabel metal1 21298 14246 21298 14246 0 _0061_
rlabel metal1 21988 14586 21988 14586 0 _0062_
rlabel metal1 22264 14790 22264 14790 0 _0063_
rlabel metal2 22264 17646 22264 17646 0 _0064_
rlabel metal1 4922 13362 4922 13362 0 _0065_
rlabel metal1 4876 17714 4876 17714 0 _0066_
rlabel metal1 19596 15470 19596 15470 0 _0067_
rlabel metal2 17066 14484 17066 14484 0 _0068_
rlabel metal1 3726 13328 3726 13328 0 _0069_
rlabel metal2 5290 20604 5290 20604 0 _0070_
rlabel metal2 5382 20638 5382 20638 0 _0071_
rlabel metal1 5152 18258 5152 18258 0 _0072_
rlabel metal1 4554 12410 4554 12410 0 _0073_
rlabel metal1 5612 22746 5612 22746 0 _0074_
rlabel metal2 6210 15878 6210 15878 0 _0075_
rlabel metal1 5704 15674 5704 15674 0 _0076_
rlabel metal1 5750 16048 5750 16048 0 _0077_
rlabel metal1 5428 22134 5428 22134 0 _0078_
rlabel metal1 7038 16082 7038 16082 0 _0079_
rlabel metal1 6532 22474 6532 22474 0 _0080_
rlabel metal1 13570 21421 13570 21421 0 _0081_
rlabel metal1 7590 21454 7590 21454 0 _0082_
rlabel metal1 8050 21590 8050 21590 0 _0083_
rlabel metal1 6900 16626 6900 16626 0 _0084_
rlabel metal1 6532 16422 6532 16422 0 _0085_
rlabel metal1 6716 16014 6716 16014 0 _0086_
rlabel metal1 6210 15912 6210 15912 0 _0087_
rlabel metal1 6210 15674 6210 15674 0 _0088_
rlabel metal1 13064 20366 13064 20366 0 _0089_
rlabel metal1 7544 15334 7544 15334 0 _0090_
rlabel metal1 6670 15674 6670 15674 0 _0091_
rlabel metal2 8786 20638 8786 20638 0 _0092_
rlabel metal1 5842 20570 5842 20570 0 _0093_
rlabel metal1 6670 18836 6670 18836 0 _0094_
rlabel metal1 7866 15436 7866 15436 0 _0095_
rlabel metal1 10166 20978 10166 20978 0 _0096_
rlabel metal1 7222 15572 7222 15572 0 _0097_
rlabel metal1 7498 14892 7498 14892 0 _0098_
rlabel metal1 7314 15130 7314 15130 0 _0099_
rlabel metal2 6762 14144 6762 14144 0 _0100_
rlabel metal1 6578 14484 6578 14484 0 _0101_
rlabel via1 7499 14453 7499 14453 0 _0102_
rlabel metal1 8786 13328 8786 13328 0 _0103_
rlabel metal1 7682 12308 7682 12308 0 _0104_
rlabel metal2 8234 15130 8234 15130 0 _0105_
rlabel metal1 14122 20978 14122 20978 0 _0106_
rlabel metal2 14674 20706 14674 20706 0 _0107_
rlabel via1 5750 19890 5750 19890 0 _0108_
rlabel metal2 7130 19516 7130 19516 0 _0109_
rlabel metal2 5842 19890 5842 19890 0 _0110_
rlabel metal1 5704 19278 5704 19278 0 _0111_
rlabel metal1 7360 19278 7360 19278 0 _0112_
rlabel metal1 9246 18836 9246 18836 0 _0113_
rlabel metal1 8970 14960 8970 14960 0 _0114_
rlabel metal1 7728 14790 7728 14790 0 _0115_
rlabel metal2 8142 14552 8142 14552 0 _0116_
rlabel metal1 7820 13906 7820 13906 0 _0117_
rlabel metal1 8602 13770 8602 13770 0 _0118_
rlabel metal1 8303 13226 8303 13226 0 _0119_
rlabel metal1 9016 13906 9016 13906 0 _0120_
rlabel metal1 8510 12410 8510 12410 0 _0121_
rlabel metal1 13340 20026 13340 20026 0 _0122_
rlabel metal1 14352 19278 14352 19278 0 _0123_
rlabel metal1 4784 19142 4784 19142 0 _0124_
rlabel metal2 6026 18054 6026 18054 0 _0125_
rlabel metal1 7038 18292 7038 18292 0 _0126_
rlabel metal1 7084 18190 7084 18190 0 _0127_
rlabel metal2 8234 17442 8234 17442 0 _0128_
rlabel metal1 9522 16694 9522 16694 0 _0129_
rlabel metal1 9476 18802 9476 18802 0 _0130_
rlabel metal1 9614 16150 9614 16150 0 _0131_
rlabel metal1 9982 15470 9982 15470 0 _0132_
rlabel metal1 10028 14450 10028 14450 0 _0133_
rlabel metal1 8510 14586 8510 14586 0 _0134_
rlabel metal1 9982 13362 9982 13362 0 _0135_
rlabel via1 10074 13770 10074 13770 0 _0136_
rlabel metal1 10396 12954 10396 12954 0 _0137_
rlabel metal1 13800 19890 13800 19890 0 _0138_
rlabel metal1 14030 19788 14030 19788 0 _0139_
rlabel metal2 6072 20978 6072 20978 0 _0140_
rlabel metal1 5888 17714 5888 17714 0 _0141_
rlabel viali 6578 18191 6578 18191 0 _0142_
rlabel metal1 8786 17748 8786 17748 0 _0143_
rlabel metal1 10258 17170 10258 17170 0 _0144_
rlabel metal2 20746 20876 20746 20876 0 _0145_
rlabel metal1 13616 18802 13616 18802 0 _0146_
rlabel metal1 7682 17714 7682 17714 0 _0147_
rlabel metal1 9614 17177 9614 17177 0 _0148_
rlabel metal1 11408 16558 11408 16558 0 _0149_
rlabel metal1 11914 14926 11914 14926 0 _0150_
rlabel metal2 11086 16048 11086 16048 0 _0151_
rlabel metal1 10856 15538 10856 15538 0 _0152_
rlabel metal1 11776 15130 11776 15130 0 _0153_
rlabel metal1 11454 14314 11454 14314 0 _0154_
rlabel metal2 12466 14246 12466 14246 0 _0155_
rlabel metal1 11362 13260 11362 13260 0 _0156_
rlabel metal1 11316 11866 11316 11866 0 _0157_
rlabel metal1 10994 16728 10994 16728 0 _0158_
rlabel metal2 11546 15844 11546 15844 0 _0159_
rlabel metal1 19688 22610 19688 22610 0 _0160_
rlabel metal1 18676 22066 18676 22066 0 _0161_
rlabel metal1 18906 22950 18906 22950 0 _0162_
rlabel metal1 9384 22610 9384 22610 0 _0163_
rlabel metal1 6394 21930 6394 21930 0 _0164_
rlabel metal1 6946 22440 6946 22440 0 _0165_
rlabel metal1 7038 22032 7038 22032 0 _0166_
rlabel metal1 6808 22066 6808 22066 0 _0167_
rlabel metal1 8004 21998 8004 21998 0 _0168_
rlabel metal1 8556 22542 8556 22542 0 _0169_
rlabel metal2 10534 22005 10534 22005 0 _0170_
rlabel metal1 10350 22202 10350 22202 0 _0171_
rlabel metal1 11224 17714 11224 17714 0 _0172_
rlabel metal2 8326 17986 8326 17986 0 _0173_
rlabel metal1 11086 17714 11086 17714 0 _0174_
rlabel metal1 11638 17170 11638 17170 0 _0175_
rlabel metal1 11684 14994 11684 14994 0 _0176_
rlabel metal2 11914 14518 11914 14518 0 _0177_
rlabel metal1 11868 13294 11868 13294 0 _0178_
rlabel metal2 12926 12818 12926 12818 0 _0179_
rlabel metal2 12466 11968 12466 11968 0 _0180_
rlabel metal1 19826 21386 19826 21386 0 _0181_
rlabel metal1 17020 22066 17020 22066 0 _0182_
rlabel metal1 16376 22950 16376 22950 0 _0183_
rlabel metal1 17664 23018 17664 23018 0 _0184_
rlabel metal1 21206 21998 21206 21998 0 _0185_
rlabel metal1 8142 21454 8142 21454 0 _0186_
rlabel metal1 8970 21658 8970 21658 0 _0187_
rlabel metal1 9522 22508 9522 22508 0 _0188_
rlabel metal1 10120 22610 10120 22610 0 _0189_
rlabel metal1 11546 22576 11546 22576 0 _0190_
rlabel metal1 10902 21998 10902 21998 0 _0191_
rlabel metal1 12466 22474 12466 22474 0 _0192_
rlabel metal1 12650 16728 12650 16728 0 _0193_
rlabel metal1 12190 17170 12190 17170 0 _0194_
rlabel metal1 14122 15028 14122 15028 0 _0195_
rlabel metal1 13616 14246 13616 14246 0 _0196_
rlabel metal1 12788 14994 12788 14994 0 _0197_
rlabel metal2 12834 14722 12834 14722 0 _0198_
rlabel metal1 13248 14450 13248 14450 0 _0199_
rlabel metal1 13984 12818 13984 12818 0 _0200_
rlabel metal1 14812 12886 14812 12886 0 _0201_
rlabel metal1 12742 22576 12742 22576 0 _0202_
rlabel via1 12633 16626 12633 16626 0 _0203_
rlabel metal1 22126 21896 22126 21896 0 _0204_
rlabel metal1 13800 19278 13800 19278 0 _0205_
rlabel metal1 12926 20400 12926 20400 0 _0206_
rlabel metal1 12880 20570 12880 20570 0 _0207_
rlabel metal1 8326 20978 8326 20978 0 _0208_
rlabel metal1 10396 20978 10396 20978 0 _0209_
rlabel metal2 10994 21182 10994 21182 0 _0210_
rlabel metal2 12742 21080 12742 21080 0 _0211_
rlabel metal1 11638 22066 11638 22066 0 _0212_
rlabel metal1 13570 21991 13570 21991 0 _0213_
rlabel metal2 12558 16898 12558 16898 0 _0214_
rlabel metal1 13156 14858 13156 14858 0 _0215_
rlabel metal1 13708 14382 13708 14382 0 _0216_
rlabel metal1 14076 13906 14076 13906 0 _0217_
rlabel metal2 14858 13192 14858 13192 0 _0218_
rlabel metal1 14076 12410 14076 12410 0 _0219_
rlabel metal1 8878 19312 8878 19312 0 _0220_
rlabel metal1 8464 18870 8464 18870 0 _0221_
rlabel metal1 9430 19278 9430 19278 0 _0222_
rlabel metal1 12834 19822 12834 19822 0 _0223_
rlabel metal1 11270 21012 11270 21012 0 _0224_
rlabel metal2 11638 20332 11638 20332 0 _0225_
rlabel metal1 13938 19278 13938 19278 0 _0226_
rlabel metal1 14076 17646 14076 17646 0 _0227_
rlabel metal1 13432 21114 13432 21114 0 _0228_
rlabel metal1 14122 17510 14122 17510 0 _0229_
rlabel metal1 15042 16490 15042 16490 0 _0230_
rlabel metal2 12466 15062 12466 15062 0 _0231_
rlabel metal1 13064 14586 13064 14586 0 _0232_
rlabel metal1 14398 16626 14398 16626 0 _0233_
rlabel metal1 14582 16150 14582 16150 0 _0234_
rlabel metal1 13478 15606 13478 15606 0 _0235_
rlabel metal1 14398 15470 14398 15470 0 _0236_
rlabel metal1 15456 13906 15456 13906 0 _0237_
rlabel metal1 15318 12750 15318 12750 0 _0238_
rlabel viali 12548 19278 12548 19278 0 _0239_
rlabel metal1 13570 18224 13570 18224 0 _0240_
rlabel metal1 11822 18802 11822 18802 0 _0241_
rlabel metal1 11178 18700 11178 18700 0 _0242_
rlabel metal1 12098 18700 12098 18700 0 _0243_
rlabel metal1 13662 17850 13662 17850 0 _0244_
rlabel metal2 15134 16796 15134 16796 0 _0245_
rlabel metal2 14766 16966 14766 16966 0 _0246_
rlabel metal2 15042 16524 15042 16524 0 _0247_
rlabel metal1 15732 12750 15732 12750 0 _0248_
rlabel metal1 16238 12954 16238 12954 0 _0249_
rlabel metal1 5198 20434 5198 20434 0 _0250_
rlabel metal2 7774 20332 7774 20332 0 _0251_
rlabel metal2 10258 19618 10258 19618 0 _0252_
rlabel metal1 13478 18768 13478 18768 0 _0253_
rlabel metal1 14674 18802 14674 18802 0 _0254_
rlabel metal1 14858 18258 14858 18258 0 _0255_
rlabel metal1 16146 18224 16146 18224 0 _0256_
rlabel metal1 16146 17170 16146 17170 0 _0257_
rlabel metal1 12006 18224 12006 18224 0 _0258_
rlabel metal1 15180 17102 15180 17102 0 _0259_
rlabel metal1 16652 16014 16652 16014 0 _0260_
rlabel metal1 14674 15980 14674 15980 0 _0261_
rlabel metal1 13386 17816 13386 17816 0 _0262_
rlabel viali 16790 17102 16790 17102 0 _0263_
rlabel metal1 16284 16014 16284 16014 0 _0264_
rlabel metal1 16974 15436 16974 15436 0 _0265_
rlabel metal1 16698 15470 16698 15470 0 _0266_
rlabel metal2 17802 15300 17802 15300 0 _0267_
rlabel metal1 17342 20944 17342 20944 0 _0268_
rlabel metal1 17526 21012 17526 21012 0 _0269_
rlabel metal1 17066 19890 17066 19890 0 _0270_
rlabel metal1 17618 19346 17618 19346 0 _0271_
rlabel metal1 11638 19244 11638 19244 0 _0272_
rlabel metal1 16974 19278 16974 19278 0 _0273_
rlabel metal1 17434 18802 17434 18802 0 _0274_
rlabel metal1 16652 16626 16652 16626 0 _0275_
rlabel metal1 15364 18258 15364 18258 0 _0276_
rlabel metal1 16836 16558 16836 16558 0 _0277_
rlabel metal1 17204 16558 17204 16558 0 _0278_
rlabel metal1 17066 17000 17066 17000 0 _0279_
rlabel metal1 16882 16082 16882 16082 0 _0280_
rlabel metal1 17572 14586 17572 14586 0 _0281_
rlabel metal1 16560 13838 16560 13838 0 _0282_
rlabel metal1 17526 19958 17526 19958 0 _0283_
rlabel metal1 17618 19958 17618 19958 0 _0284_
rlabel metal1 16790 22406 16790 22406 0 _0285_
rlabel metal1 18860 21998 18860 21998 0 _0286_
rlabel metal1 17710 22134 17710 22134 0 _0287_
rlabel metal1 17802 21522 17802 21522 0 _0288_
rlabel metal1 18078 21522 18078 21522 0 _0289_
rlabel metal1 18492 20366 18492 20366 0 _0290_
rlabel metal1 18906 19856 18906 19856 0 _0291_
rlabel metal1 18446 19890 18446 19890 0 _0292_
rlabel metal1 18722 19346 18722 19346 0 _0293_
rlabel metal1 19734 18836 19734 18836 0 _0294_
rlabel metal1 17940 18870 17940 18870 0 _0295_
rlabel metal1 19435 18802 19435 18802 0 _0296_
rlabel metal1 18722 17748 18722 17748 0 _0297_
rlabel metal1 16882 16422 16882 16422 0 _0298_
rlabel metal1 18308 17034 18308 17034 0 _0299_
rlabel metal1 17273 17102 17273 17102 0 _0300_
rlabel metal1 16698 17170 16698 17170 0 _0301_
rlabel metal1 18170 17000 18170 17000 0 _0302_
rlabel metal1 18998 17238 18998 17238 0 _0303_
rlabel metal2 20102 16320 20102 16320 0 _0304_
rlabel metal1 18354 15028 18354 15028 0 _0305_
rlabel metal1 19642 19958 19642 19958 0 _0306_
rlabel metal1 21206 22950 21206 22950 0 _0307_
rlabel metal1 20240 23154 20240 23154 0 _0308_
rlabel metal2 19596 21692 19596 21692 0 _0309_
rlabel metal1 19964 21658 19964 21658 0 _0310_
rlabel metal1 20332 22066 20332 22066 0 _0311_
rlabel metal1 19596 21522 19596 21522 0 _0312_
rlabel metal2 18722 20740 18722 20740 0 _0313_
rlabel metal2 18768 19210 18768 19210 0 _0314_
rlabel metal1 19320 19414 19320 19414 0 _0315_
rlabel metal1 18998 17748 18998 17748 0 _0316_
rlabel metal1 18814 17680 18814 17680 0 _0317_
rlabel metal1 19550 18700 19550 18700 0 _0318_
rlabel metal1 18998 16592 18998 16592 0 _0319_
rlabel metal1 18998 15674 18998 15674 0 _0320_
rlabel metal1 19964 14926 19964 14926 0 _0321_
rlabel metal2 20654 18054 20654 18054 0 _0322_
rlabel metal2 20378 19108 20378 19108 0 _0323_
rlabel metal1 19550 21114 19550 21114 0 _0324_
rlabel metal1 22402 21522 22402 21522 0 _0325_
rlabel metal1 21390 22610 21390 22610 0 _0326_
rlabel metal1 22494 21930 22494 21930 0 _0327_
rlabel metal1 21896 22066 21896 22066 0 _0328_
rlabel metal1 22356 22202 22356 22202 0 _0329_
rlabel metal2 22126 21964 22126 21964 0 _0330_
rlabel metal1 22402 20434 22402 20434 0 _0331_
rlabel metal2 22586 20842 22586 20842 0 _0332_
rlabel metal1 22287 20298 22287 20298 0 _0333_
rlabel metal1 22494 19278 22494 19278 0 _0334_
rlabel metal1 20516 18258 20516 18258 0 _0335_
rlabel metal1 20654 17850 20654 17850 0 _0336_
rlabel metal2 22218 19448 22218 19448 0 _0337_
rlabel metal1 21344 19890 21344 19890 0 _0338_
rlabel metal1 21482 21012 21482 21012 0 _0339_
rlabel metal1 21068 20978 21068 20978 0 _0340_
rlabel viali 22130 20366 22130 20366 0 _0341_
rlabel metal1 20884 20366 20884 20366 0 _0342_
rlabel metal2 22310 19754 22310 19754 0 _0343_
rlabel via1 21873 18394 21873 18394 0 _0344_
rlabel metal2 22126 18768 22126 18768 0 _0345_
rlabel metal1 22218 18224 22218 18224 0 _0346_
rlabel metal1 21298 19346 21298 19346 0 _0347_
rlabel metal1 21298 19482 21298 19482 0 _0348_
rlabel metal2 20838 19754 20838 19754 0 _0349_
rlabel metal1 21298 19244 21298 19244 0 _0350_
rlabel metal1 20930 17714 20930 17714 0 _0351_
rlabel metal1 21482 18088 21482 18088 0 _0352_
rlabel metal2 21390 17442 21390 17442 0 _0353_
rlabel metal1 21436 17850 21436 17850 0 _0354_
rlabel metal1 5980 10030 5980 10030 0 _0355_
rlabel metal1 6578 10234 6578 10234 0 _0356_
rlabel metal1 5980 10982 5980 10982 0 _0357_
rlabel metal1 6072 11186 6072 11186 0 _0358_
rlabel metal1 6256 10982 6256 10982 0 _0359_
rlabel metal2 6578 10812 6578 10812 0 _0360_
rlabel metal2 5566 10812 5566 10812 0 _0361_
rlabel metal1 6164 10506 6164 10506 0 _0362_
rlabel metal1 9338 10608 9338 10608 0 _0363_
rlabel metal1 7092 11322 7092 11322 0 _0364_
rlabel metal1 8050 10608 8050 10608 0 _0365_
rlabel metal1 7820 10574 7820 10574 0 _0366_
rlabel metal1 8648 10778 8648 10778 0 _0367_
rlabel metal2 8694 11084 8694 11084 0 _0368_
rlabel metal2 9890 10812 9890 10812 0 _0369_
rlabel metal1 9430 10030 9430 10030 0 _0370_
rlabel metal1 9246 10540 9246 10540 0 _0371_
rlabel metal1 8326 10132 8326 10132 0 _0372_
rlabel metal1 8924 10234 8924 10234 0 _0373_
rlabel metal1 12052 9486 12052 9486 0 _0374_
rlabel metal1 9614 10642 9614 10642 0 _0375_
rlabel metal1 9982 10030 9982 10030 0 _0376_
rlabel metal2 10626 9792 10626 9792 0 _0377_
rlabel metal1 10580 10642 10580 10642 0 _0378_
rlabel metal1 11224 10098 11224 10098 0 _0379_
rlabel metal1 11362 9554 11362 9554 0 _0380_
rlabel metal1 12190 9588 12190 9588 0 _0381_
rlabel metal1 10994 9554 10994 9554 0 _0382_
rlabel metal1 12098 9384 12098 9384 0 _0383_
rlabel metal1 13524 9622 13524 9622 0 _0384_
rlabel metal2 12650 10880 12650 10880 0 _0385_
rlabel metal1 13248 9554 13248 9554 0 _0386_
rlabel metal1 14168 9690 14168 9690 0 _0387_
rlabel metal1 14168 10642 14168 10642 0 _0388_
rlabel metal1 14720 10574 14720 10574 0 _0389_
rlabel metal1 14766 9554 14766 9554 0 _0390_
rlabel metal2 14306 9860 14306 9860 0 _0391_
rlabel metal2 13938 9690 13938 9690 0 _0392_
rlabel metal1 14168 9146 14168 9146 0 _0393_
rlabel metal1 16376 10234 16376 10234 0 _0394_
rlabel metal1 16146 11220 16146 11220 0 _0395_
rlabel metal1 16192 10642 16192 10642 0 _0396_
rlabel metal1 17112 10778 17112 10778 0 _0397_
rlabel metal1 16422 11764 16422 11764 0 _0398_
rlabel metal1 16882 11186 16882 11186 0 _0399_
rlabel metal2 16790 10812 16790 10812 0 _0400_
rlabel metal1 17894 10676 17894 10676 0 _0401_
rlabel metal1 17066 10642 17066 10642 0 _0402_
rlabel metal1 17756 10506 17756 10506 0 _0403_
rlabel metal1 19274 10778 19274 10778 0 _0404_
rlabel metal1 18170 12308 18170 12308 0 _0405_
rlabel metal1 18538 11730 18538 11730 0 _0406_
rlabel metal1 19642 11866 19642 11866 0 _0407_
rlabel metal1 19366 12818 19366 12818 0 _0408_
rlabel metal1 20102 11764 20102 11764 0 _0409_
rlabel metal1 20010 13396 20010 13396 0 _0410_
rlabel metal2 20102 12789 20102 12789 0 _0411_
rlabel metal1 19642 11118 19642 11118 0 _0412_
rlabel metal1 20700 11866 20700 11866 0 _0413_
rlabel metal1 21101 13498 21101 13498 0 _0414_
rlabel metal2 21298 12614 21298 12614 0 _0415_
rlabel metal1 21206 12206 21206 12206 0 _0416_
rlabel metal1 21436 12818 21436 12818 0 _0417_
rlabel metal1 21206 12342 21206 12342 0 _0418_
rlabel metal1 22034 12240 22034 12240 0 _0419_
rlabel metal1 22402 14484 22402 14484 0 _0420_
rlabel metal1 22356 12818 22356 12818 0 _0421_
rlabel metal1 21942 12886 21942 12886 0 _0422_
rlabel metal1 21850 14280 21850 14280 0 _0423_
rlabel metal1 22310 12614 22310 12614 0 _0424_
rlabel metal2 22126 6392 22126 6392 0 _0425_
rlabel metal1 21206 6358 21206 6358 0 _0426_
rlabel metal2 22586 7106 22586 7106 0 _0427_
rlabel metal1 21206 6834 21206 6834 0 _0428_
rlabel metal1 21712 6970 21712 6970 0 _0429_
rlabel metal1 22172 7514 22172 7514 0 _0430_
rlabel metal1 21896 12410 21896 12410 0 _0431_
rlabel metal1 20976 11322 20976 11322 0 _0432_
rlabel metal1 20562 8908 20562 8908 0 _0433_
rlabel metal1 4830 5168 4830 5168 0 _0434_
rlabel metal1 6716 4658 6716 4658 0 _0435_
rlabel metal1 6302 5814 6302 5814 0 _0436_
rlabel metal1 14490 7956 14490 7956 0 _0437_
rlabel metal1 7209 5882 7209 5882 0 _0438_
rlabel metal1 7038 5610 7038 5610 0 _0439_
rlabel metal1 5566 6766 5566 6766 0 _0440_
rlabel metal1 4968 6834 4968 6834 0 _0441_
rlabel metal1 4922 8466 4922 8466 0 _0442_
rlabel metal1 5842 8602 5842 8602 0 _0443_
rlabel metal2 6578 9792 6578 9792 0 _0444_
rlabel metal1 4186 9486 4186 9486 0 _0445_
rlabel metal2 6486 8874 6486 8874 0 _0446_
rlabel metal1 20286 9520 20286 9520 0 _0447_
rlabel metal1 6302 8364 6302 8364 0 _0448_
rlabel metal1 7360 8330 7360 8330 0 _0449_
rlabel metal1 8234 7412 8234 7412 0 _0450_
rlabel metal1 8050 7514 8050 7514 0 _0451_
rlabel metal1 7544 7310 7544 7310 0 _0452_
rlabel via1 10810 8466 10810 8466 0 _0453_
rlabel metal1 8786 7276 8786 7276 0 _0454_
rlabel metal1 9798 7242 9798 7242 0 _0455_
rlabel metal1 9890 7820 9890 7820 0 _0456_
rlabel metal1 10074 7514 10074 7514 0 _0457_
rlabel metal1 10488 6834 10488 6834 0 _0458_
rlabel metal1 11546 7344 11546 7344 0 _0459_
rlabel metal1 11684 7310 11684 7310 0 _0460_
rlabel metal1 12696 7514 12696 7514 0 _0461_
rlabel metal2 14858 7650 14858 7650 0 _0462_
rlabel metal1 14950 7718 14950 7718 0 _0463_
rlabel metal1 14306 7854 14306 7854 0 _0464_
rlabel metal1 14076 8534 14076 8534 0 _0465_
rlabel metal1 14444 6834 14444 6834 0 _0466_
rlabel metal1 16928 7990 16928 7990 0 _0467_
rlabel metal1 16652 8534 16652 8534 0 _0468_
rlabel metal1 15732 8602 15732 8602 0 _0469_
rlabel metal1 15916 6834 15916 6834 0 _0470_
rlabel metal1 16744 9486 16744 9486 0 _0471_
rlabel metal2 17710 9010 17710 9010 0 _0472_
rlabel metal1 19044 9010 19044 9010 0 _0473_
rlabel metal1 19320 9622 19320 9622 0 _0474_
rlabel metal1 20010 8806 20010 8806 0 _0475_
rlabel metal1 19182 9146 19182 9146 0 _0476_
rlabel metal2 19734 9894 19734 9894 0 _0477_
rlabel metal1 20056 9690 20056 9690 0 _0478_
rlabel metal1 20884 10234 20884 10234 0 _0479_
rlabel metal1 20654 9622 20654 9622 0 _0480_
rlabel metal1 21068 10778 21068 10778 0 _0481_
rlabel metal2 22126 10948 22126 10948 0 _0482_
rlabel metal1 21712 9894 21712 9894 0 _0483_
rlabel metal1 21206 9520 21206 9520 0 _0484_
rlabel metal1 20608 8398 20608 8398 0 _0485_
rlabel metal1 22034 8296 22034 8296 0 _0486_
rlabel metal1 21252 8602 21252 8602 0 _0487_
rlabel metal1 22494 8466 22494 8466 0 _0488_
rlabel metal1 19228 6834 19228 6834 0 _0489_
rlabel metal1 21804 5134 21804 5134 0 _0490_
rlabel metal1 18768 6630 18768 6630 0 _0491_
rlabel metal2 18170 5780 18170 5780 0 _0492_
rlabel metal1 18308 6834 18308 6834 0 _0493_
rlabel metal1 18354 6222 18354 6222 0 _0494_
rlabel metal1 18078 6256 18078 6256 0 _0495_
rlabel metal2 19918 7123 19918 7123 0 _0496_
rlabel metal1 20608 6426 20608 6426 0 _0497_
rlabel metal1 20470 4726 20470 4726 0 _0498_
rlabel metal1 20654 6256 20654 6256 0 _0499_
rlabel metal1 21436 14926 21436 14926 0 _0500_
rlabel metal2 23046 3961 23046 3961 0 clk_in
rlabel metal1 22540 18938 22540 18938 0 clk_out
rlabel metal1 6394 6154 6394 6154 0 count\[0\]
rlabel metal2 10534 9248 10534 9248 0 count\[10\]
rlabel metal1 11040 8262 11040 8262 0 count\[11\]
rlabel metal1 11040 8398 11040 8398 0 count\[12\]
rlabel metal1 13662 8534 13662 8534 0 count\[13\]
rlabel metal2 14214 8772 14214 8772 0 count\[14\]
rlabel metal1 14950 8330 14950 8330 0 count\[15\]
rlabel metal1 16192 8466 16192 8466 0 count\[16\]
rlabel metal1 16514 8432 16514 8432 0 count\[17\]
rlabel metal1 17434 9146 17434 9146 0 count\[18\]
rlabel metal2 18814 10540 18814 10540 0 count\[19\]
rlabel metal1 4692 6222 4692 6222 0 count\[1\]
rlabel metal1 19642 9486 19642 9486 0 count\[20\]
rlabel metal1 19090 9520 19090 9520 0 count\[21\]
rlabel metal1 21114 12750 21114 12750 0 count\[22\]
rlabel metal1 21252 11866 21252 11866 0 count\[23\]
rlabel metal1 21942 12750 21942 12750 0 count\[24\]
rlabel metal1 22448 10098 22448 10098 0 count\[25\]
rlabel metal1 21666 8058 21666 8058 0 count\[26\]
rlabel metal2 22586 6052 22586 6052 0 count\[27\]
rlabel metal1 18998 6834 18998 6834 0 count\[28\]
rlabel metal1 19642 6800 19642 6800 0 count\[29\]
rlabel metal1 5980 6766 5980 6766 0 count\[2\]
rlabel metal2 21390 5780 21390 5780 0 count\[30\]
rlabel metal1 20286 6834 20286 6834 0 count\[31\]
rlabel metal1 6348 6426 6348 6426 0 count\[3\]
rlabel metal1 6256 10030 6256 10030 0 count\[4\]
rlabel metal2 5750 10370 5750 10370 0 count\[5\]
rlabel metal1 6164 9486 6164 9486 0 count\[6\]
rlabel via1 7774 10523 7774 10523 0 count\[7\]
rlabel metal2 8602 9248 8602 9248 0 count\[8\]
rlabel metal1 8694 8432 8694 8432 0 count\[9\]
rlabel metal1 13202 8942 13202 8942 0 net1
rlabel metal1 19826 22066 19826 22066 0 net10
rlabel metal1 14214 15538 14214 15538 0 net11
rlabel metal1 15364 20366 15364 20366 0 net12
rlabel metal1 20700 22542 20700 22542 0 net13
rlabel metal1 5290 19142 5290 19142 0 net14
rlabel metal1 10626 12716 10626 12716 0 net15
rlabel metal1 22448 18190 22448 18190 0 net16
rlabel metal1 4324 9010 4324 9010 0 net17
rlabel metal1 13984 7310 13984 7310 0 net18
rlabel metal1 13938 8806 13938 8806 0 net19
rlabel metal1 14490 12648 14490 12648 0 net2
rlabel metal2 19642 10540 19642 10540 0 net20
rlabel via2 21298 9044 21298 9044 0 net21
rlabel metal1 23000 16218 23000 16218 0 net22
rlabel metal1 22678 7310 22678 7310 0 net23
rlabel metal1 5060 22066 5060 22066 0 net3
rlabel metal1 4324 19822 4324 19822 0 net4
rlabel metal1 15916 20978 15916 20978 0 net5
rlabel metal2 14490 21216 14490 21216 0 net6
rlabel metal1 20286 22508 20286 22508 0 net7
rlabel metal1 20792 21386 20792 21386 0 net8
rlabel metal1 20976 21658 20976 21658 0 net9
rlabel metal1 23184 12274 23184 12274 0 nrst
rlabel metal1 1748 23154 1748 23154 0 scale[0]
rlabel metal1 4738 23222 4738 23222 0 scale[1]
rlabel metal1 7682 23222 7682 23222 0 scale[2]
rlabel metal1 10856 23222 10856 23222 0 scale[3]
rlabel metal1 13524 23154 13524 23154 0 scale[4]
rlabel metal1 17710 23188 17710 23188 0 scale[5]
rlabel metal2 19458 23443 19458 23443 0 scale[6]
rlabel metal1 22356 23154 22356 23154 0 scale[7]
rlabel metal2 22034 15130 22034 15130 0 signal_clk_out
rlabel metal1 7866 12206 7866 12206 0 true_scale\[10\]
rlabel metal1 8464 12614 8464 12614 0 true_scale\[11\]
rlabel metal1 10902 11186 10902 11186 0 true_scale\[12\]
rlabel metal1 11086 11730 11086 11730 0 true_scale\[13\]
rlabel metal2 12374 11832 12374 11832 0 true_scale\[14\]
rlabel metal1 13754 11866 13754 11866 0 true_scale\[15\]
rlabel metal1 14950 12750 14950 12750 0 true_scale\[16\]
rlabel metal1 15778 13702 15778 13702 0 true_scale\[17\]
rlabel metal2 17618 12954 17618 12954 0 true_scale\[18\]
rlabel metal1 17894 14790 17894 14790 0 true_scale\[19\]
rlabel metal1 17986 14042 17986 14042 0 true_scale\[20\]
rlabel metal1 20056 15130 20056 15130 0 true_scale\[21\]
rlabel metal2 18446 15062 18446 15062 0 true_scale\[22\]
rlabel metal1 20838 16966 20838 16966 0 true_scale\[23\]
rlabel metal1 21758 17850 21758 17850 0 true_scale\[24\]
rlabel metal1 22816 17238 22816 17238 0 true_scale\[25\]
rlabel metal2 22678 17544 22678 17544 0 true_scale\[26\]
rlabel metal1 5980 13498 5980 13498 0 true_scale\[5\]
rlabel metal1 5428 14450 5428 14450 0 true_scale\[6\]
rlabel via1 5566 12342 5566 12342 0 true_scale\[7\]
rlabel metal1 5842 15334 5842 15334 0 true_scale\[8\]
rlabel metal1 6394 15130 6394 15130 0 true_scale\[9\]
flabel metal4 3760 23760 3800 23820 0 FreeSans 320 90 0 0 VPWR
flabel metal4 19130 23510 19160 23580 0 FreeSans 320 90 0 0 VGND
<< properties >>
string FIXED_BBOX 0 0 24000 24000
<< end >>
