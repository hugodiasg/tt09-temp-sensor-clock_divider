magic
tech sky130A
magscale 1 2
timestamp 1729283362
<< viali >>
rect 7665 23273 7699 23307
rect 11069 23205 11103 23239
rect 18705 23205 18739 23239
rect 18905 23205 18939 23239
rect 19717 23205 19751 23239
rect 20637 23205 20671 23239
rect 20853 23205 20887 23239
rect 1777 23137 1811 23171
rect 5089 23137 5123 23171
rect 5181 23137 5215 23171
rect 5825 23137 5859 23171
rect 6009 23137 6043 23171
rect 6469 23137 6503 23171
rect 6561 23137 6595 23171
rect 6745 23137 6779 23171
rect 7849 23137 7883 23171
rect 8677 23137 8711 23171
rect 8861 23137 8895 23171
rect 13553 23137 13587 23171
rect 16497 23137 16531 23171
rect 19165 23137 19199 23171
rect 19349 23137 19383 23171
rect 19441 23137 19475 23171
rect 21281 23137 21315 23171
rect 21465 23137 21499 23171
rect 22385 23137 22419 23171
rect 6285 23069 6319 23103
rect 13737 23069 13771 23103
rect 22569 23069 22603 23103
rect 1961 23001 1995 23035
rect 6653 23001 6687 23035
rect 9045 23001 9079 23035
rect 4905 22933 4939 22967
rect 5365 22933 5399 22967
rect 11345 22933 11379 22967
rect 16681 22933 16715 22967
rect 18889 22933 18923 22967
rect 19073 22933 19107 22967
rect 19165 22933 19199 22967
rect 20821 22933 20855 22967
rect 21005 22933 21039 22967
rect 21649 22933 21683 22967
rect 8033 22729 8067 22763
rect 9781 22729 9815 22763
rect 12541 22729 12575 22763
rect 12817 22729 12851 22763
rect 15485 22729 15519 22763
rect 17693 22729 17727 22763
rect 20453 22729 20487 22763
rect 21557 22729 21591 22763
rect 4721 22661 4755 22695
rect 7757 22661 7791 22695
rect 10149 22661 10183 22695
rect 11253 22661 11287 22695
rect 15669 22661 15703 22695
rect 18429 22661 18463 22695
rect 21097 22661 21131 22695
rect 22017 22661 22051 22695
rect 5273 22593 5307 22627
rect 9137 22593 9171 22627
rect 10333 22593 10367 22627
rect 14013 22593 14047 22627
rect 16221 22593 16255 22627
rect 17417 22593 17451 22627
rect 17969 22593 18003 22627
rect 18521 22593 18555 22627
rect 19165 22593 19199 22627
rect 20821 22593 20855 22627
rect 21557 22593 21591 22627
rect 21741 22593 21775 22627
rect 4629 22525 4663 22559
rect 4905 22525 4939 22559
rect 5917 22525 5951 22559
rect 6377 22525 6411 22559
rect 7481 22525 7515 22559
rect 7573 22525 7607 22559
rect 7757 22525 7791 22559
rect 8493 22525 8527 22559
rect 8677 22525 8711 22559
rect 8769 22525 8803 22559
rect 8861 22525 8895 22559
rect 9229 22525 9263 22559
rect 9321 22525 9355 22559
rect 9505 22525 9539 22559
rect 9597 22525 9631 22559
rect 10517 22525 10551 22559
rect 10610 22525 10644 22559
rect 10977 22525 11011 22559
rect 12817 22525 12851 22559
rect 12909 22525 12943 22559
rect 13553 22525 13587 22559
rect 13646 22525 13680 22559
rect 14197 22525 14231 22559
rect 17049 22525 17083 22559
rect 18153 22525 18187 22559
rect 18981 22525 19015 22559
rect 19809 22525 19843 22559
rect 20177 22525 20211 22559
rect 20269 22525 20303 22559
rect 20453 22525 20487 22559
rect 20729 22525 20763 22559
rect 21189 22525 21223 22559
rect 21281 22525 21315 22559
rect 21465 22525 21499 22559
rect 7849 22457 7883 22491
rect 9873 22457 9907 22491
rect 11253 22457 11287 22491
rect 12357 22457 12391 22491
rect 15301 22457 15335 22491
rect 16957 22457 16991 22491
rect 17233 22457 17267 22491
rect 17509 22457 17543 22491
rect 8054 22389 8088 22423
rect 8217 22389 8251 22423
rect 10885 22389 10919 22423
rect 11069 22389 11103 22423
rect 12557 22389 12591 22423
rect 12725 22389 12759 22423
rect 13185 22389 13219 22423
rect 13921 22389 13955 22423
rect 14381 22389 14415 22423
rect 15511 22389 15545 22423
rect 17709 22389 17743 22423
rect 17877 22389 17911 22423
rect 22201 22389 22235 22423
rect 4813 22185 4847 22219
rect 5273 22185 5307 22219
rect 9229 22185 9263 22219
rect 12541 22185 12575 22219
rect 14565 22185 14599 22219
rect 15301 22185 15335 22219
rect 4629 22117 4663 22151
rect 5365 22117 5399 22151
rect 19993 22117 20027 22151
rect 21833 22117 21867 22151
rect 22477 22117 22511 22151
rect 22661 22117 22695 22151
rect 6837 22049 6871 22083
rect 7205 22049 7239 22083
rect 8125 22049 8159 22083
rect 8953 22049 8987 22083
rect 9781 22049 9815 22083
rect 9965 22049 9999 22083
rect 10793 22049 10827 22083
rect 12081 22049 12115 22083
rect 12633 22049 12667 22083
rect 13001 22049 13035 22083
rect 14933 22049 14967 22083
rect 15761 22049 15795 22083
rect 16129 22049 16163 22083
rect 16773 22049 16807 22083
rect 17049 22049 17083 22083
rect 17877 22049 17911 22083
rect 18521 22049 18555 22083
rect 19257 22049 19291 22083
rect 19901 22049 19935 22083
rect 20177 22049 20211 22083
rect 20453 22049 20487 22083
rect 21925 22049 21959 22083
rect 22109 22049 22143 22083
rect 22201 22049 22235 22083
rect 22385 22049 22419 22083
rect 8033 21981 8067 22015
rect 9045 21981 9079 22015
rect 9413 21981 9447 22015
rect 11253 21981 11287 22015
rect 12173 21981 12207 22015
rect 12357 21981 12391 22015
rect 13277 21981 13311 22015
rect 13829 21981 13863 22015
rect 14105 21981 14139 22015
rect 14197 21981 14231 22015
rect 15025 21981 15059 22015
rect 15669 21981 15703 22015
rect 17969 21981 18003 22015
rect 20361 21981 20395 22015
rect 21741 21981 21775 22015
rect 22293 21981 22327 22015
rect 7113 21913 7147 21947
rect 15393 21913 15427 21947
rect 21465 21913 21499 21947
rect 22385 21913 22419 21947
rect 4813 21845 4847 21879
rect 4997 21845 5031 21879
rect 9413 21845 9447 21879
rect 13921 21845 13955 21879
rect 16313 21845 16347 21879
rect 17601 21845 17635 21879
rect 18705 21845 18739 21879
rect 19809 21845 19843 21879
rect 20545 21845 20579 21879
rect 21281 21845 21315 21879
rect 12265 21641 12299 21675
rect 12541 21641 12575 21675
rect 16681 21641 16715 21675
rect 9137 21573 9171 21607
rect 12449 21573 12483 21607
rect 16221 21573 16255 21607
rect 17509 21573 17543 21607
rect 18245 21573 18279 21607
rect 21465 21573 21499 21607
rect 10885 21505 10919 21539
rect 12357 21505 12391 21539
rect 13185 21505 13219 21539
rect 14381 21505 14415 21539
rect 15025 21505 15059 21539
rect 15209 21505 15243 21539
rect 15761 21505 15795 21539
rect 17601 21505 17635 21539
rect 18061 21505 18095 21539
rect 18797 21505 18831 21539
rect 21741 21505 21775 21539
rect 5273 21437 5307 21471
rect 6745 21437 6779 21471
rect 7297 21437 7331 21471
rect 7665 21437 7699 21471
rect 7757 21437 7791 21471
rect 7941 21437 7975 21471
rect 8033 21437 8067 21471
rect 8493 21437 8527 21471
rect 8677 21437 8711 21471
rect 8953 21437 8987 21471
rect 9229 21437 9263 21471
rect 9321 21437 9355 21471
rect 9597 21437 9631 21471
rect 9965 21437 9999 21471
rect 10149 21437 10183 21471
rect 10333 21437 10367 21471
rect 10517 21437 10551 21471
rect 10701 21437 10735 21471
rect 10977 21437 11011 21471
rect 11437 21437 11471 21471
rect 11713 21437 11747 21471
rect 11989 21437 12023 21471
rect 12081 21437 12115 21471
rect 12265 21437 12299 21471
rect 12633 21437 12667 21471
rect 13093 21437 13127 21471
rect 14197 21437 14231 21471
rect 14933 21437 14967 21471
rect 15117 21437 15151 21471
rect 15853 21437 15887 21471
rect 16313 21437 16347 21471
rect 16497 21437 16531 21471
rect 16957 21437 16991 21471
rect 17141 21437 17175 21471
rect 17233 21437 17267 21471
rect 17325 21437 17359 21471
rect 17509 21437 17543 21471
rect 17969 21437 18003 21471
rect 18521 21437 18555 21471
rect 18705 21437 18739 21471
rect 20360 21437 20394 21471
rect 20453 21437 20487 21471
rect 20545 21437 20579 21471
rect 20638 21437 20672 21471
rect 21005 21437 21039 21471
rect 21189 21437 21223 21471
rect 4537 21369 4571 21403
rect 8217 21369 8251 21403
rect 9781 21369 9815 21403
rect 10609 21369 10643 21403
rect 11529 21369 11563 21403
rect 15393 21369 15427 21403
rect 15577 21369 15611 21403
rect 18245 21369 18279 21403
rect 21097 21369 21131 21403
rect 9413 21301 9447 21335
rect 11345 21301 11379 21335
rect 11897 21301 11931 21335
rect 12725 21301 12759 21335
rect 13369 21301 13403 21335
rect 13553 21301 13587 21335
rect 16773 21301 16807 21335
rect 18429 21301 18463 21335
rect 20085 21301 20119 21335
rect 20913 21301 20947 21335
rect 21281 21301 21315 21335
rect 6929 21097 6963 21131
rect 8217 21097 8251 21131
rect 10425 21097 10459 21131
rect 15761 21097 15795 21131
rect 16681 21097 16715 21131
rect 18061 21097 18095 21131
rect 20897 21097 20931 21131
rect 16221 21029 16255 21063
rect 17693 21029 17727 21063
rect 20637 21029 20671 21063
rect 21097 21029 21131 21063
rect 5457 20961 5491 20995
rect 5641 20961 5675 20995
rect 6009 20961 6043 20995
rect 7389 20961 7423 20995
rect 7481 20961 7515 20995
rect 7665 20961 7699 20995
rect 8401 20961 8435 20995
rect 9137 20961 9171 20995
rect 9321 20961 9355 20995
rect 9413 20961 9447 20995
rect 9505 20961 9539 20995
rect 9689 20961 9723 20995
rect 10057 20961 10091 20995
rect 10241 20961 10275 20995
rect 10333 20961 10367 20995
rect 10517 20961 10551 20995
rect 15669 20961 15703 20995
rect 15945 20961 15979 20995
rect 16129 20961 16163 20995
rect 16313 20961 16347 20995
rect 16497 20961 16531 20995
rect 16681 20961 16715 20995
rect 17877 20961 17911 20995
rect 20085 20961 20119 20995
rect 20269 20961 20303 20995
rect 20361 20961 20395 20995
rect 20453 20961 20487 20995
rect 21465 20961 21499 20995
rect 21649 20961 21683 20995
rect 21741 20961 21775 20995
rect 6101 20893 6135 20927
rect 7021 20893 7055 20927
rect 7205 20893 7239 20927
rect 8493 20893 8527 20927
rect 8861 20893 8895 20927
rect 13553 20893 13587 20927
rect 14289 20893 14323 20927
rect 21557 20893 21591 20927
rect 15945 20825 15979 20859
rect 5549 20757 5583 20791
rect 6377 20757 6411 20791
rect 6561 20757 6595 20791
rect 7849 20757 7883 20791
rect 8953 20757 8987 20791
rect 9597 20757 9631 20791
rect 10057 20757 10091 20791
rect 20177 20757 20211 20791
rect 20637 20757 20671 20791
rect 20729 20757 20763 20791
rect 20913 20757 20947 20791
rect 21281 20757 21315 20791
rect 6837 20553 6871 20587
rect 20637 20553 20671 20587
rect 5089 20485 5123 20519
rect 10701 20485 10735 20519
rect 10241 20417 10275 20451
rect 11805 20417 11839 20451
rect 21005 20417 21039 20451
rect 4445 20349 4479 20383
rect 4629 20349 4663 20383
rect 4721 20349 4755 20383
rect 4813 20349 4847 20383
rect 4905 20349 4939 20383
rect 5457 20349 5491 20383
rect 5641 20349 5675 20383
rect 5825 20349 5859 20383
rect 5917 20349 5951 20383
rect 6101 20349 6135 20383
rect 6745 20349 6779 20383
rect 10333 20349 10367 20383
rect 11989 20349 12023 20383
rect 12633 20349 12667 20383
rect 12725 20349 12759 20383
rect 19441 20349 19475 20383
rect 19533 20349 19567 20383
rect 20545 20349 20579 20383
rect 20637 20349 20671 20383
rect 21373 20349 21407 20383
rect 21465 20349 21499 20383
rect 21649 20349 21683 20383
rect 19257 20281 19291 20315
rect 21833 20281 21867 20315
rect 22477 20281 22511 20315
rect 4261 20213 4295 20247
rect 6009 20213 6043 20247
rect 12173 20213 12207 20247
rect 12909 20213 12943 20247
rect 19533 20213 19567 20247
rect 20913 20213 20947 20247
rect 21925 20213 21959 20247
rect 22385 20213 22419 20247
rect 5089 20009 5123 20043
rect 21465 20009 21499 20043
rect 4077 19941 4111 19975
rect 4629 19941 4663 19975
rect 17325 19941 17359 19975
rect 17601 19941 17635 19975
rect 17801 19941 17835 19975
rect 19073 19941 19107 19975
rect 5181 19873 5215 19907
rect 5273 19873 5307 19907
rect 6009 19873 6043 19907
rect 7021 19873 7055 19907
rect 10333 19873 10367 19907
rect 10701 19873 10735 19907
rect 11989 19873 12023 19907
rect 12449 19873 12483 19907
rect 13185 19873 13219 19907
rect 13645 19873 13679 19907
rect 13783 19873 13817 19907
rect 16497 19873 16531 19907
rect 16957 19873 16991 19907
rect 17050 19873 17084 19907
rect 18337 19873 18371 19907
rect 18429 19873 18463 19907
rect 18981 19873 19015 19907
rect 19257 19873 19291 19907
rect 19717 19873 19751 19907
rect 20177 19873 20211 19907
rect 20545 19873 20579 19907
rect 20821 19873 20855 19907
rect 21005 19873 21039 19907
rect 21462 19873 21496 19907
rect 22293 19873 22327 19907
rect 22385 19873 22419 19907
rect 22569 19873 22603 19907
rect 4537 19805 4571 19839
rect 6101 19805 6135 19839
rect 6745 19805 6779 19839
rect 8861 19805 8895 19839
rect 13093 19805 13127 19839
rect 16405 19805 16439 19839
rect 18153 19805 18187 19839
rect 18245 19805 18279 19839
rect 18613 19805 18647 19839
rect 19441 19805 19475 19839
rect 19809 19805 19843 19839
rect 19901 19805 19935 19839
rect 19993 19805 20027 19839
rect 20637 19805 20671 19839
rect 21925 19805 21959 19839
rect 23029 19805 23063 19839
rect 4353 19737 4387 19771
rect 4905 19737 4939 19771
rect 6377 19737 6411 19771
rect 6837 19737 6871 19771
rect 7205 19737 7239 19771
rect 13553 19737 13587 19771
rect 16865 19737 16899 19771
rect 5181 19669 5215 19703
rect 5549 19669 5583 19703
rect 13829 19669 13863 19703
rect 17785 19669 17819 19703
rect 17969 19669 18003 19703
rect 19533 19669 19567 19703
rect 20361 19669 20395 19703
rect 21281 19669 21315 19703
rect 21833 19669 21867 19703
rect 4537 19465 4571 19499
rect 5273 19465 5307 19499
rect 9689 19465 9723 19499
rect 11989 19465 12023 19499
rect 13369 19465 13403 19499
rect 14381 19465 14415 19499
rect 18705 19465 18739 19499
rect 22201 19465 22235 19499
rect 7573 19397 7607 19431
rect 12173 19397 12207 19431
rect 12725 19397 12759 19431
rect 13001 19397 13035 19431
rect 14933 19397 14967 19431
rect 18153 19397 18187 19431
rect 4169 19329 4203 19363
rect 4721 19329 4755 19363
rect 5181 19329 5215 19363
rect 5365 19329 5399 19363
rect 7113 19329 7147 19363
rect 11713 19329 11747 19363
rect 12541 19329 12575 19363
rect 12909 19329 12943 19363
rect 13645 19329 13679 19363
rect 14105 19329 14139 19363
rect 14289 19329 14323 19363
rect 16865 19329 16899 19363
rect 17325 19329 17359 19363
rect 4261 19261 4295 19295
rect 4353 19261 4387 19295
rect 4813 19261 4847 19295
rect 5273 19261 5307 19295
rect 6285 19261 6319 19295
rect 6469 19261 6503 19295
rect 7205 19261 7239 19295
rect 7665 19261 7699 19295
rect 7849 19261 7883 19295
rect 8033 19261 8067 19295
rect 8769 19261 8803 19295
rect 8861 19261 8895 19295
rect 9045 19261 9079 19295
rect 10241 19261 10275 19295
rect 10977 19261 11011 19295
rect 11621 19261 11655 19295
rect 12081 19261 12115 19295
rect 12265 19261 12299 19295
rect 12817 19261 12851 19295
rect 13185 19261 13219 19295
rect 13737 19261 13771 19295
rect 14197 19261 14231 19295
rect 14657 19261 14691 19295
rect 14933 19261 14967 19295
rect 16773 19261 16807 19295
rect 17233 19261 17267 19295
rect 17417 19261 17451 19295
rect 17877 19261 17911 19295
rect 17969 19261 18003 19295
rect 18153 19261 18187 19295
rect 18245 19261 18279 19295
rect 18429 19261 18463 19295
rect 18705 19261 18739 19295
rect 18889 19261 18923 19295
rect 19165 19261 19199 19295
rect 20821 19261 20855 19295
rect 21088 19261 21122 19295
rect 22477 19261 22511 19295
rect 22661 19261 22695 19295
rect 22845 19261 22879 19295
rect 6101 19193 6135 19227
rect 7941 19193 7975 19227
rect 8401 19193 8435 19227
rect 14749 19193 14783 19227
rect 19432 19193 19466 19227
rect 22569 19193 22603 19227
rect 5641 19125 5675 19159
rect 8217 19125 8251 19159
rect 12817 19125 12851 19159
rect 14565 19125 14599 19159
rect 17141 19125 17175 19159
rect 18337 19125 18371 19159
rect 20545 19125 20579 19159
rect 22293 19125 22327 19159
rect 7481 18921 7515 18955
rect 7941 18921 7975 18955
rect 12725 18921 12759 18955
rect 13369 18921 13403 18955
rect 18061 18921 18095 18955
rect 19993 18921 20027 18955
rect 20637 18921 20671 18955
rect 22753 18921 22787 18955
rect 5273 18853 5307 18887
rect 9597 18853 9631 18887
rect 16221 18853 16255 18887
rect 21640 18853 21674 18887
rect 5181 18785 5215 18819
rect 5457 18785 5491 18819
rect 6653 18785 6687 18819
rect 7573 18785 7607 18819
rect 7757 18785 7791 18819
rect 8493 18785 8527 18819
rect 8953 18785 8987 18819
rect 9413 18785 9447 18819
rect 10057 18785 10091 18819
rect 10425 18785 10459 18819
rect 11345 18785 11379 18819
rect 11805 18785 11839 18819
rect 12357 18785 12391 18819
rect 13093 18785 13127 18819
rect 13737 18785 13771 18819
rect 14289 18785 14323 18819
rect 14933 18785 14967 18819
rect 15761 18785 15795 18819
rect 16129 18785 16163 18819
rect 16405 18785 16439 18819
rect 17693 18785 17727 18819
rect 17785 18785 17819 18819
rect 17969 18785 18003 18819
rect 18153 18785 18187 18819
rect 20177 18785 20211 18819
rect 20361 18785 20395 18819
rect 20545 18785 20579 18819
rect 21097 18785 21131 18819
rect 23029 18785 23063 18819
rect 6561 18717 6595 18751
rect 8585 18717 8619 18751
rect 8861 18717 8895 18751
rect 10333 18717 10367 18751
rect 11069 18717 11103 18751
rect 12265 18717 12299 18751
rect 13185 18717 13219 18751
rect 13369 18717 13403 18751
rect 14013 18717 14047 18751
rect 14197 18717 14231 18751
rect 14841 18717 14875 18751
rect 15301 18717 15335 18751
rect 15853 18717 15887 18751
rect 21373 18717 21407 18751
rect 5457 18649 5491 18683
rect 8125 18649 8159 18683
rect 9321 18649 9355 18683
rect 9965 18649 9999 18683
rect 10793 18649 10827 18683
rect 11805 18649 11839 18683
rect 13553 18649 13587 18683
rect 16405 18649 16439 18683
rect 20913 18649 20947 18683
rect 9781 18581 9815 18615
rect 13921 18581 13955 18615
rect 14565 18581 14599 18615
rect 15485 18581 15519 18615
rect 17509 18581 17543 18615
rect 22937 18581 22971 18615
rect 5365 18377 5399 18411
rect 7113 18377 7147 18411
rect 14933 18377 14967 18411
rect 15577 18377 15611 18411
rect 17785 18377 17819 18411
rect 18061 18377 18095 18411
rect 21557 18377 21591 18411
rect 23029 18377 23063 18411
rect 4629 18309 4663 18343
rect 17601 18309 17635 18343
rect 18981 18309 19015 18343
rect 5549 18241 5583 18275
rect 6193 18241 6227 18275
rect 11713 18241 11747 18275
rect 11989 18241 12023 18275
rect 14381 18241 14415 18275
rect 14657 18241 14691 18275
rect 15209 18241 15243 18275
rect 17969 18241 18003 18275
rect 18429 18241 18463 18275
rect 18889 18241 18923 18275
rect 4077 18173 4111 18207
rect 4445 18173 4479 18207
rect 4721 18173 4755 18207
rect 4905 18173 4939 18207
rect 5181 18173 5215 18207
rect 5641 18173 5675 18207
rect 6101 18173 6135 18207
rect 6285 18173 6319 18207
rect 6653 18173 6687 18207
rect 6929 18173 6963 18207
rect 8585 18173 8619 18207
rect 8769 18173 8803 18207
rect 8861 18173 8895 18207
rect 9045 18173 9079 18207
rect 10793 18173 10827 18207
rect 10977 18173 11011 18207
rect 11161 18173 11195 18207
rect 11253 18173 11287 18207
rect 11897 18173 11931 18207
rect 14289 18173 14323 18207
rect 14749 18173 14783 18207
rect 14933 18173 14967 18207
rect 15393 18173 15427 18207
rect 17417 18173 17451 18207
rect 17601 18173 17635 18207
rect 17693 18173 17727 18207
rect 18245 18173 18279 18207
rect 18797 18173 18831 18207
rect 19073 18173 19107 18207
rect 19257 18173 19291 18207
rect 19349 18173 19383 18207
rect 19717 18173 19751 18207
rect 21281 18173 21315 18207
rect 21649 18173 21683 18207
rect 4261 18105 4295 18139
rect 4353 18105 4387 18139
rect 6745 18105 6779 18139
rect 11437 18105 11471 18139
rect 17969 18105 18003 18139
rect 19533 18105 19567 18139
rect 19625 18105 19659 18139
rect 21557 18105 21591 18139
rect 21916 18105 21950 18139
rect 6009 18037 6043 18071
rect 8769 18037 8803 18071
rect 8861 18037 8895 18071
rect 19901 18037 19935 18071
rect 21373 18037 21407 18071
rect 4077 17833 4111 17867
rect 9137 17833 9171 17867
rect 10057 17833 10091 17867
rect 18245 17833 18279 17867
rect 18613 17833 18647 17867
rect 22753 17833 22787 17867
rect 3801 17765 3835 17799
rect 19748 17765 19782 17799
rect 21097 17765 21131 17799
rect 21526 17765 21560 17799
rect 4353 17697 4387 17731
rect 4629 17697 4663 17731
rect 5181 17697 5215 17731
rect 5917 17697 5951 17731
rect 6101 17697 6135 17731
rect 6929 17697 6963 17731
rect 7389 17697 7423 17731
rect 7573 17697 7607 17731
rect 9045 17697 9079 17731
rect 9321 17697 9355 17731
rect 9689 17697 9723 17731
rect 16313 17697 16347 17731
rect 16497 17697 16531 17731
rect 16589 17697 16623 17731
rect 17233 17697 17267 17731
rect 17417 17697 17451 17731
rect 17601 17697 17635 17731
rect 17877 17697 17911 17731
rect 18153 17697 18187 17731
rect 18337 17697 18371 17731
rect 18521 17697 18555 17731
rect 19993 17697 20027 17731
rect 20913 17697 20947 17731
rect 22937 17697 22971 17731
rect 23029 17697 23063 17731
rect 4445 17629 4479 17663
rect 4997 17629 5031 17663
rect 5549 17629 5583 17663
rect 9781 17629 9815 17663
rect 20637 17629 20671 17663
rect 21281 17629 21315 17663
rect 22753 17629 22787 17663
rect 5457 17561 5491 17595
rect 4721 17493 4755 17527
rect 7573 17493 7607 17527
rect 9321 17493 9355 17527
rect 16129 17493 16163 17527
rect 16681 17493 16715 17527
rect 18337 17493 18371 17527
rect 20729 17493 20763 17527
rect 22661 17493 22695 17527
rect 4537 17289 4571 17323
rect 5457 17289 5491 17323
rect 5641 17289 5675 17323
rect 9505 17289 9539 17323
rect 13921 17289 13955 17323
rect 15945 17289 15979 17323
rect 17141 17289 17175 17323
rect 17509 17289 17543 17323
rect 18337 17289 18371 17323
rect 22385 17289 22419 17323
rect 4997 17221 5031 17255
rect 12541 17221 12575 17255
rect 13369 17221 13403 17255
rect 16865 17221 16899 17255
rect 5181 17153 5215 17187
rect 6009 17153 6043 17187
rect 6285 17153 6319 17187
rect 7297 17153 7331 17187
rect 8217 17153 8251 17187
rect 9689 17153 9723 17187
rect 10149 17153 10183 17187
rect 10609 17153 10643 17187
rect 11805 17153 11839 17187
rect 12081 17153 12115 17187
rect 12909 17153 12943 17187
rect 14933 17153 14967 17187
rect 15761 17153 15795 17187
rect 18199 17153 18233 17187
rect 4169 17085 4203 17119
rect 4629 17085 4663 17119
rect 4997 17085 5031 17119
rect 5917 17085 5951 17119
rect 7389 17085 7423 17119
rect 8861 17085 8895 17119
rect 9137 17085 9171 17119
rect 9321 17085 9355 17119
rect 9781 17085 9815 17119
rect 10241 17085 10275 17119
rect 10701 17085 10735 17119
rect 10885 17085 10919 17119
rect 11713 17085 11747 17119
rect 12173 17085 12207 17119
rect 13001 17085 13035 17119
rect 13737 17085 13771 17119
rect 15025 17085 15059 17119
rect 16037 17085 16071 17119
rect 16313 17085 16347 17119
rect 16589 17085 16623 17119
rect 16773 17085 16807 17119
rect 16865 17085 16899 17119
rect 17049 17085 17083 17119
rect 17141 17085 17175 17119
rect 17233 17085 17267 17119
rect 18061 17085 18095 17119
rect 18521 17085 18555 17119
rect 18705 17085 18739 17119
rect 4353 17017 4387 17051
rect 5273 17017 5307 17051
rect 10793 17017 10827 17051
rect 11161 17017 11195 17051
rect 13553 17017 13587 17051
rect 16129 17017 16163 17051
rect 18429 17017 18463 17051
rect 18950 17017 18984 17051
rect 22661 17017 22695 17051
rect 5473 16949 5507 16983
rect 8677 16949 8711 16983
rect 11713 16949 11747 16983
rect 15393 16949 15427 16983
rect 15485 16949 15519 16983
rect 20085 16949 20119 16983
rect 4261 16745 4295 16779
rect 9045 16745 9079 16779
rect 9613 16745 9647 16779
rect 14565 16745 14599 16779
rect 16497 16745 16531 16779
rect 18889 16745 18923 16779
rect 4879 16677 4913 16711
rect 4997 16677 5031 16711
rect 5549 16677 5583 16711
rect 9413 16677 9447 16711
rect 13185 16677 13219 16711
rect 14105 16677 14139 16711
rect 14749 16677 14783 16711
rect 15117 16677 15151 16711
rect 16129 16677 16163 16711
rect 16345 16677 16379 16711
rect 16681 16677 16715 16711
rect 21833 16677 21867 16711
rect 4169 16609 4203 16643
rect 5089 16609 5123 16643
rect 5181 16609 5215 16643
rect 5457 16609 5491 16643
rect 7481 16609 7515 16643
rect 8861 16609 8895 16643
rect 9137 16609 9171 16643
rect 9321 16609 9355 16643
rect 13093 16609 13127 16643
rect 13277 16609 13311 16643
rect 13369 16609 13403 16643
rect 13553 16609 13587 16643
rect 13645 16609 13679 16643
rect 13737 16609 13771 16643
rect 13921 16609 13955 16643
rect 14289 16609 14323 16643
rect 14381 16609 14415 16643
rect 14657 16609 14691 16643
rect 15025 16609 15059 16643
rect 15209 16609 15243 16643
rect 16589 16609 16623 16643
rect 18797 16609 18831 16643
rect 18981 16609 19015 16643
rect 21557 16609 21591 16643
rect 4629 16541 4663 16575
rect 4721 16541 4755 16575
rect 7389 16541 7423 16575
rect 13461 16541 13495 16575
rect 15301 16541 15335 16575
rect 15485 16541 15519 16575
rect 21833 16541 21867 16575
rect 4445 16473 4479 16507
rect 7849 16473 7883 16507
rect 14933 16473 14967 16507
rect 5365 16405 5399 16439
rect 9597 16405 9631 16439
rect 9781 16405 9815 16439
rect 15393 16405 15427 16439
rect 16313 16405 16347 16439
rect 21649 16405 21683 16439
rect 13369 16201 13403 16235
rect 19165 16201 19199 16235
rect 21833 16201 21867 16235
rect 22569 16201 22603 16235
rect 6929 16133 6963 16167
rect 12541 16133 12575 16167
rect 14473 16133 14507 16167
rect 15393 16133 15427 16167
rect 16957 16133 16991 16167
rect 19809 16133 19843 16167
rect 5365 16065 5399 16099
rect 5641 16065 5675 16099
rect 6653 16065 6687 16099
rect 6837 16065 6871 16099
rect 11253 16065 11287 16099
rect 11713 16065 11747 16099
rect 13645 16065 13679 16099
rect 15301 16065 15335 16099
rect 16313 16065 16347 16099
rect 16405 16065 16439 16099
rect 19625 16065 19659 16099
rect 21281 16065 21315 16099
rect 21557 16065 21591 16099
rect 21741 16065 21775 16099
rect 5273 15997 5307 16031
rect 5733 15997 5767 16031
rect 5917 15997 5951 16031
rect 6561 15997 6595 16031
rect 7113 15997 7147 16031
rect 7205 15997 7239 16031
rect 11345 15997 11379 16031
rect 11805 15997 11839 16031
rect 11989 15997 12023 16031
rect 12265 15997 12299 16031
rect 13185 15997 13219 16031
rect 13737 15997 13771 16031
rect 14197 15997 14231 16031
rect 14473 15997 14507 16031
rect 15209 15997 15243 16031
rect 15485 15997 15519 16031
rect 16129 15997 16163 16031
rect 16221 15997 16255 16031
rect 16681 15997 16715 16031
rect 16773 15997 16807 16031
rect 16957 15997 16991 16031
rect 19165 15997 19199 16031
rect 19257 15997 19291 16031
rect 19901 15997 19935 16031
rect 20269 15997 20303 16031
rect 20545 15997 20579 16031
rect 20729 15997 20763 16031
rect 21189 15997 21223 16031
rect 21649 15997 21683 16031
rect 22385 15997 22419 16031
rect 6929 15929 6963 15963
rect 12173 15929 12207 15963
rect 12541 15929 12575 15963
rect 13001 15929 13035 15963
rect 15669 15929 15703 15963
rect 20085 15929 20119 15963
rect 22201 15929 22235 15963
rect 5917 15861 5951 15895
rect 6193 15861 6227 15895
rect 12357 15861 12391 15895
rect 14105 15861 14139 15895
rect 14289 15861 14323 15895
rect 16589 15861 16623 15895
rect 19533 15861 19567 15895
rect 19625 15861 19659 15895
rect 20453 15861 20487 15895
rect 20729 15861 20763 15895
rect 22017 15861 22051 15895
rect 4445 15657 4479 15691
rect 20821 15657 20855 15691
rect 16497 15589 16531 15623
rect 20269 15589 20303 15623
rect 20485 15589 20519 15623
rect 4077 15521 4111 15555
rect 4261 15521 4295 15555
rect 5273 15521 5307 15555
rect 6009 15521 6043 15555
rect 6653 15521 6687 15555
rect 7297 15521 7331 15555
rect 8861 15521 8895 15555
rect 9321 15521 9355 15555
rect 9414 15521 9448 15555
rect 9965 15521 9999 15555
rect 10058 15521 10092 15555
rect 11713 15521 11747 15555
rect 13001 15521 13035 15555
rect 13369 15521 13403 15555
rect 16313 15521 16347 15555
rect 16405 15521 16439 15555
rect 16681 15521 16715 15555
rect 16957 15521 16991 15555
rect 17049 15521 17083 15555
rect 17325 15521 17359 15555
rect 19533 15521 19567 15555
rect 19717 15521 19751 15555
rect 20729 15521 20763 15555
rect 21005 15521 21039 15555
rect 21741 15521 21775 15555
rect 5181 15453 5215 15487
rect 6101 15453 6135 15487
rect 6745 15453 6779 15487
rect 7205 15453 7239 15487
rect 8769 15453 8803 15487
rect 11621 15453 11655 15487
rect 13921 15453 13955 15487
rect 21649 15453 21683 15487
rect 5641 15385 5675 15419
rect 6377 15385 6411 15419
rect 7021 15385 7055 15419
rect 7665 15385 7699 15419
rect 9229 15385 9263 15419
rect 12081 15385 12115 15419
rect 9505 15317 9539 15351
rect 10149 15317 10183 15351
rect 16129 15317 16163 15351
rect 16773 15317 16807 15351
rect 17233 15317 17267 15351
rect 19625 15317 19659 15351
rect 20453 15317 20487 15351
rect 20637 15317 20671 15351
rect 21005 15317 21039 15351
rect 22109 15317 22143 15351
rect 6561 15113 6595 15147
rect 12725 15113 12759 15147
rect 14105 15113 14139 15147
rect 17049 15113 17083 15147
rect 18245 15113 18279 15147
rect 20545 15113 20579 15147
rect 5089 15045 5123 15079
rect 6377 15045 6411 15079
rect 7941 15045 7975 15079
rect 20729 15045 20763 15079
rect 21741 15045 21775 15079
rect 22017 15045 22051 15079
rect 6101 14977 6135 15011
rect 7481 14977 7515 15011
rect 9689 14977 9723 15011
rect 10517 14977 10551 15011
rect 11437 14977 11471 15011
rect 17877 14977 17911 15011
rect 18705 14977 18739 15011
rect 19165 14977 19199 15011
rect 19717 14977 19751 15011
rect 19993 14977 20027 15011
rect 20361 14977 20395 15011
rect 21465 14977 21499 15011
rect 21833 14977 21867 15011
rect 22385 14977 22419 15011
rect 4629 14909 4663 14943
rect 4813 14909 4847 14943
rect 4997 14909 5031 14943
rect 5273 14909 5307 14943
rect 5365 14909 5399 14943
rect 6929 14909 6963 14943
rect 7022 14909 7056 14943
rect 7573 14909 7607 14943
rect 9781 14909 9815 14943
rect 10609 14909 10643 14943
rect 11345 14909 11379 14943
rect 11529 14909 11563 14943
rect 11989 14909 12023 14943
rect 12265 14909 12299 14943
rect 13553 14909 13587 14943
rect 13645 14909 13679 14943
rect 13829 14909 13863 14943
rect 13921 14909 13955 14943
rect 15669 14909 15703 14943
rect 15936 14909 15970 14943
rect 17693 14909 17727 14943
rect 17969 14909 18003 14943
rect 18061 14909 18095 14943
rect 19073 14909 19107 14943
rect 19625 14909 19659 14943
rect 20545 14909 20579 14943
rect 21373 14909 21407 14943
rect 21925 14909 21959 14943
rect 22293 14909 22327 14943
rect 22569 14909 22603 14943
rect 22661 14909 22695 14943
rect 4721 14841 4755 14875
rect 5089 14841 5123 14875
rect 7297 14841 7331 14875
rect 12541 14841 12575 14875
rect 12741 14841 12775 14875
rect 17509 14841 17543 14875
rect 18245 14841 18279 14875
rect 20269 14841 20303 14875
rect 22201 14841 22235 14875
rect 4445 14773 4479 14807
rect 9413 14773 9447 14807
rect 10241 14773 10275 14807
rect 12081 14773 12115 14807
rect 12449 14773 12483 14807
rect 12909 14773 12943 14807
rect 22385 14773 22419 14807
rect 10149 14569 10183 14603
rect 11069 14569 11103 14603
rect 13001 14569 13035 14603
rect 13645 14569 13679 14603
rect 17509 14569 17543 14603
rect 17693 14569 17727 14603
rect 18077 14569 18111 14603
rect 19441 14569 19475 14603
rect 23029 14569 23063 14603
rect 4506 14501 4540 14535
rect 9597 14501 9631 14535
rect 10333 14501 10367 14535
rect 10577 14501 10611 14535
rect 10767 14501 10801 14535
rect 13829 14501 13863 14535
rect 16396 14501 16430 14535
rect 17877 14501 17911 14535
rect 21649 14501 21683 14535
rect 7849 14433 7883 14467
rect 8309 14433 8343 14467
rect 8402 14433 8436 14467
rect 9137 14433 9171 14467
rect 9321 14433 9355 14467
rect 9781 14433 9815 14467
rect 10057 14433 10091 14467
rect 10977 14433 11011 14467
rect 11253 14433 11287 14467
rect 12909 14433 12943 14467
rect 13185 14433 13219 14467
rect 13369 14433 13403 14467
rect 13737 14433 13771 14467
rect 14013 14433 14047 14467
rect 17601 14433 17635 14467
rect 17785 14433 17819 14467
rect 18521 14433 18555 14467
rect 18981 14433 19015 14467
rect 19257 14433 19291 14467
rect 21281 14433 21315 14467
rect 21373 14433 21407 14467
rect 21557 14433 21591 14467
rect 21833 14433 21867 14467
rect 21925 14433 21959 14467
rect 22017 14433 22051 14467
rect 22155 14433 22189 14467
rect 22385 14433 22419 14467
rect 22845 14433 22879 14467
rect 4261 14365 4295 14399
rect 7941 14365 7975 14399
rect 13277 14365 13311 14399
rect 16129 14365 16163 14399
rect 18613 14365 18647 14399
rect 19073 14365 19107 14399
rect 22293 14365 22327 14399
rect 22661 14365 22695 14399
rect 8677 14297 8711 14331
rect 10333 14297 10367 14331
rect 18889 14297 18923 14331
rect 21557 14297 21591 14331
rect 5641 14229 5675 14263
rect 8217 14229 8251 14263
rect 9229 14229 9263 14263
rect 9965 14229 9999 14263
rect 10425 14229 10459 14263
rect 10587 14229 10621 14263
rect 11437 14229 11471 14263
rect 14197 14229 14231 14263
rect 18061 14229 18095 14263
rect 18245 14229 18279 14263
rect 19073 14229 19107 14263
rect 22477 14229 22511 14263
rect 4169 14025 4203 14059
rect 9597 14025 9631 14059
rect 10885 14025 10919 14059
rect 13829 14025 13863 14059
rect 14197 14025 14231 14059
rect 17417 14025 17451 14059
rect 17601 14025 17635 14059
rect 19073 14025 19107 14059
rect 5641 13957 5675 13991
rect 8585 13957 8619 13991
rect 9873 13957 9907 13991
rect 11069 13957 11103 13991
rect 12173 13957 12207 13991
rect 13369 13957 13403 13991
rect 14013 13957 14047 13991
rect 14289 13957 14323 13991
rect 17969 13957 18003 13991
rect 6101 13889 6135 13923
rect 6285 13889 6319 13923
rect 11161 13889 11195 13923
rect 12357 13889 12391 13923
rect 12633 13889 12667 13923
rect 12725 13889 12759 13923
rect 12817 13889 12851 13923
rect 14381 13889 14415 13923
rect 15393 13889 15427 13923
rect 20361 13889 20395 13923
rect 22201 13889 22235 13923
rect 5293 13821 5327 13855
rect 5549 13821 5583 13855
rect 8401 13821 8435 13855
rect 8585 13821 8619 13855
rect 9137 13821 9171 13855
rect 9505 13821 9539 13855
rect 9689 13821 9723 13855
rect 9965 13821 9999 13855
rect 10057 13821 10091 13855
rect 10333 13821 10367 13855
rect 10425 13821 10459 13855
rect 11345 13821 11379 13855
rect 11437 13821 11471 13855
rect 12081 13821 12115 13855
rect 12265 13821 12299 13855
rect 12541 13821 12575 13855
rect 13093 13821 13127 13855
rect 13369 13821 13403 13855
rect 14105 13821 14139 13855
rect 15577 13821 15611 13855
rect 17693 13821 17727 13855
rect 17785 13821 17819 13855
rect 17969 13821 18003 13855
rect 18889 13821 18923 13855
rect 20628 13821 20662 13855
rect 22017 13821 22051 13855
rect 10931 13787 10965 13821
rect 13875 13787 13909 13821
rect 6009 13753 6043 13787
rect 8953 13753 8987 13787
rect 9229 13753 9263 13787
rect 10241 13753 10275 13787
rect 10701 13753 10735 13787
rect 13645 13753 13679 13787
rect 15669 13753 15703 13787
rect 17233 13753 17267 13787
rect 18705 13753 18739 13787
rect 8769 13685 8803 13719
rect 10609 13685 10643 13719
rect 11161 13685 11195 13719
rect 13185 13685 13219 13719
rect 16037 13685 16071 13719
rect 17433 13685 17467 13719
rect 21741 13685 21775 13719
rect 21833 13685 21867 13719
rect 5365 13481 5399 13515
rect 6285 13481 6319 13515
rect 8309 13481 8343 13515
rect 10425 13481 10459 13515
rect 12449 13481 12483 13515
rect 12817 13481 12851 13515
rect 14565 13481 14599 13515
rect 16773 13481 16807 13515
rect 17141 13481 17175 13515
rect 18153 13481 18187 13515
rect 22385 13481 22419 13515
rect 8125 13413 8159 13447
rect 8769 13413 8803 13447
rect 15700 13413 15734 13447
rect 17969 13413 18003 13447
rect 18245 13413 18279 13447
rect 18445 13413 18479 13447
rect 19809 13413 19843 13447
rect 21557 13413 21591 13447
rect 22477 13413 22511 13447
rect 5273 13345 5307 13379
rect 6193 13345 6227 13379
rect 8401 13345 8435 13379
rect 8953 13345 8987 13379
rect 9229 13345 9263 13379
rect 9413 13345 9447 13379
rect 9965 13345 9999 13379
rect 10149 13345 10183 13379
rect 10241 13345 10275 13379
rect 10425 13345 10459 13379
rect 12357 13345 12391 13379
rect 12633 13345 12667 13379
rect 13093 13345 13127 13379
rect 13247 13345 13281 13379
rect 13829 13345 13863 13379
rect 13921 13345 13955 13379
rect 16405 13345 16439 13379
rect 16865 13345 16899 13379
rect 17785 13345 17819 13379
rect 20361 13345 20395 13379
rect 21741 13345 21775 13379
rect 22017 13345 22051 13379
rect 22201 13345 22235 13379
rect 22661 13345 22695 13379
rect 5549 13277 5583 13311
rect 6377 13277 6411 13311
rect 13461 13277 13495 13311
rect 13737 13277 13771 13311
rect 14013 13277 14047 13311
rect 15945 13277 15979 13311
rect 16497 13277 16531 13311
rect 16957 13277 16991 13311
rect 17141 13277 17175 13311
rect 20453 13277 20487 13311
rect 20545 13277 20579 13311
rect 20637 13277 20671 13311
rect 18613 13209 18647 13243
rect 20177 13209 20211 13243
rect 22845 13209 22879 13243
rect 4905 13141 4939 13175
rect 5825 13141 5859 13175
rect 8125 13141 8159 13175
rect 9137 13141 9171 13175
rect 9321 13141 9355 13175
rect 9781 13141 9815 13175
rect 13553 13141 13587 13175
rect 16589 13141 16623 13175
rect 18429 13141 18463 13175
rect 19625 13141 19659 13175
rect 19809 13141 19843 13175
rect 20821 13141 20855 13175
rect 21925 13141 21959 13175
rect 5917 12937 5951 12971
rect 12449 12937 12483 12971
rect 18061 12937 18095 12971
rect 18705 12937 18739 12971
rect 20821 12937 20855 12971
rect 20913 12937 20947 12971
rect 21097 12937 21131 12971
rect 21741 12937 21775 12971
rect 21465 12869 21499 12903
rect 21925 12869 21959 12903
rect 8677 12801 8711 12835
rect 9229 12801 9263 12835
rect 11161 12801 11195 12835
rect 11253 12801 11287 12835
rect 22017 12801 22051 12835
rect 4537 12733 4571 12767
rect 4804 12733 4838 12767
rect 6009 12733 6043 12767
rect 8585 12733 8619 12767
rect 8861 12733 8895 12767
rect 9137 12733 9171 12767
rect 9321 12733 9355 12767
rect 11345 12733 11379 12767
rect 11437 12733 11471 12767
rect 11989 12733 12023 12767
rect 12541 12733 12575 12767
rect 13553 12733 13587 12767
rect 13809 12733 13843 12767
rect 18429 12733 18463 12767
rect 18889 12733 18923 12767
rect 19165 12733 19199 12767
rect 19441 12733 19475 12767
rect 19708 12733 19742 12767
rect 22293 12733 22327 12767
rect 6276 12665 6310 12699
rect 9045 12665 9079 12699
rect 12081 12665 12115 12699
rect 18061 12665 18095 12699
rect 21557 12665 21591 12699
rect 7389 12597 7423 12631
rect 10977 12597 11011 12631
rect 12265 12597 12299 12631
rect 14933 12597 14967 12631
rect 17877 12597 17911 12631
rect 19073 12597 19107 12631
rect 21097 12597 21131 12631
rect 21757 12597 21791 12631
rect 5641 12393 5675 12427
rect 6469 12393 6503 12427
rect 6929 12393 6963 12427
rect 11345 12393 11379 12427
rect 13185 12393 13219 12427
rect 14105 12393 14139 12427
rect 15209 12393 15243 12427
rect 17601 12393 17635 12427
rect 19073 12393 19107 12427
rect 20545 12393 20579 12427
rect 21005 12393 21039 12427
rect 21649 12393 21683 12427
rect 4528 12325 4562 12359
rect 6837 12325 6871 12359
rect 8033 12325 8067 12359
rect 8401 12325 8435 12359
rect 12072 12325 12106 12359
rect 17233 12325 17267 12359
rect 17449 12325 17483 12359
rect 17960 12325 17994 12359
rect 19410 12325 19444 12359
rect 21373 12325 21407 12359
rect 4261 12257 4295 12291
rect 8125 12257 8159 12291
rect 8217 12257 8251 12291
rect 8493 12257 8527 12291
rect 8585 12257 8619 12291
rect 9229 12257 9263 12291
rect 9781 12257 9815 12291
rect 11526 12257 11560 12291
rect 11805 12257 11839 12291
rect 14289 12257 14323 12291
rect 14473 12257 14507 12291
rect 15117 12257 15151 12291
rect 16313 12257 16347 12291
rect 16957 12257 16991 12291
rect 17141 12257 17175 12291
rect 20821 12257 20855 12291
rect 22762 12257 22796 12291
rect 7021 12189 7055 12223
rect 9137 12189 9171 12223
rect 9689 12189 9723 12223
rect 11713 12189 11747 12223
rect 15301 12189 15335 12223
rect 16405 12189 16439 12223
rect 17693 12189 17727 12223
rect 19165 12189 19199 12223
rect 20637 12189 20671 12223
rect 23029 12189 23063 12223
rect 10149 12121 10183 12155
rect 8769 12053 8803 12087
rect 8953 12053 8987 12087
rect 14749 12053 14783 12087
rect 16681 12053 16715 12087
rect 17049 12053 17083 12087
rect 17417 12053 17451 12087
rect 21465 12053 21499 12087
rect 5641 11849 5675 11883
rect 9781 11849 9815 11883
rect 12081 11849 12115 11883
rect 14197 11849 14231 11883
rect 15761 11849 15795 11883
rect 17877 11849 17911 11883
rect 19717 11849 19751 11883
rect 21281 11849 21315 11883
rect 5549 11781 5583 11815
rect 5457 11713 5491 11747
rect 21557 11713 21591 11747
rect 5733 11645 5767 11679
rect 8401 11645 8435 11679
rect 8668 11645 8702 11679
rect 10701 11645 10735 11679
rect 10968 11645 11002 11679
rect 14013 11645 14047 11679
rect 14289 11645 14323 11679
rect 14381 11645 14415 11679
rect 14648 11645 14682 11679
rect 18061 11645 18095 11679
rect 19901 11645 19935 11679
rect 20545 11645 20579 11679
rect 20637 11645 20671 11679
rect 20821 11645 20855 11679
rect 20913 11645 20947 11679
rect 18245 11577 18279 11611
rect 20085 11577 20119 11611
rect 20361 11577 20395 11611
rect 21802 11577 21836 11611
rect 13829 11509 13863 11543
rect 20177 11509 20211 11543
rect 20729 11509 20763 11543
rect 21281 11509 21315 11543
rect 21465 11509 21499 11543
rect 22937 11509 22971 11543
rect 7849 11305 7883 11339
rect 14841 11305 14875 11339
rect 17877 11305 17911 11339
rect 20821 11305 20855 11339
rect 22017 11305 22051 11339
rect 22267 11305 22301 11339
rect 5917 11237 5951 11271
rect 13728 11237 13762 11271
rect 17201 11237 17235 11271
rect 17417 11237 17451 11271
rect 21833 11237 21867 11271
rect 22477 11237 22511 11271
rect 5089 11169 5123 11203
rect 6193 11169 6227 11203
rect 8033 11169 8067 11203
rect 8125 11169 8159 11203
rect 8392 11169 8426 11203
rect 10977 11169 11011 11203
rect 11244 11169 11278 11203
rect 13461 11169 13495 11203
rect 14933 11169 14967 11203
rect 15117 11169 15151 11203
rect 15209 11169 15243 11203
rect 16589 11169 16623 11203
rect 17509 11169 17543 11203
rect 19441 11169 19475 11203
rect 19708 11169 19742 11203
rect 21465 11169 21499 11203
rect 22753 11169 22787 11203
rect 5181 11101 5215 11135
rect 6009 11101 6043 11135
rect 16681 11101 16715 11135
rect 22569 11101 22603 11135
rect 5457 11033 5491 11067
rect 6377 11033 6411 11067
rect 15393 11033 15427 11067
rect 5917 10965 5951 10999
rect 9505 10965 9539 10999
rect 12357 10965 12391 10999
rect 14933 10965 14967 10999
rect 16865 10965 16899 10999
rect 17049 10965 17083 10999
rect 17233 10965 17267 10999
rect 17877 10965 17911 10999
rect 18061 10965 18095 10999
rect 21833 10965 21867 10999
rect 22109 10965 22143 10999
rect 22293 10965 22327 10999
rect 5365 10761 5399 10795
rect 5641 10761 5675 10795
rect 5825 10761 5859 10795
rect 6561 10761 6595 10795
rect 7113 10761 7147 10795
rect 8677 10761 8711 10795
rect 9597 10761 9631 10795
rect 9965 10761 9999 10795
rect 11345 10761 11379 10795
rect 11667 10761 11701 10795
rect 12081 10761 12115 10795
rect 12541 10761 12575 10795
rect 14795 10761 14829 10795
rect 16865 10761 16899 10795
rect 17141 10761 17175 10795
rect 19809 10761 19843 10795
rect 19993 10761 20027 10795
rect 21557 10761 21591 10795
rect 22845 10761 22879 10795
rect 5549 10693 5583 10727
rect 6745 10693 6779 10727
rect 11805 10693 11839 10727
rect 16497 10693 16531 10727
rect 21373 10693 21407 10727
rect 9137 10625 9171 10659
rect 9321 10625 9355 10659
rect 9597 10625 9631 10659
rect 10793 10625 10827 10659
rect 10885 10625 10919 10659
rect 12173 10625 12207 10659
rect 14933 10625 14967 10659
rect 15025 10625 15059 10659
rect 16681 10625 16715 10659
rect 18521 10625 18555 10659
rect 5825 10557 5859 10591
rect 6009 10557 6043 10591
rect 6377 10557 6411 10591
rect 6561 10557 6595 10591
rect 6837 10557 6871 10591
rect 6929 10557 6963 10591
rect 7205 10557 7239 10591
rect 7389 10557 7423 10591
rect 9045 10557 9079 10591
rect 9781 10557 9815 10591
rect 10977 10557 11011 10591
rect 11529 10557 11563 10591
rect 11989 10557 12023 10591
rect 12357 10557 12391 10591
rect 12725 10557 12759 10591
rect 12909 10557 12943 10591
rect 13093 10557 13127 10591
rect 13277 10557 13311 10591
rect 13921 10557 13955 10591
rect 14105 10557 14139 10591
rect 14289 10557 14323 10591
rect 14381 10557 14415 10591
rect 14657 10557 14691 10591
rect 15117 10557 15151 10591
rect 16221 10557 16255 10591
rect 16313 10557 16347 10591
rect 16497 10557 16531 10591
rect 16865 10557 16899 10591
rect 18254 10557 18288 10591
rect 23029 10557 23063 10591
rect 5181 10489 5215 10523
rect 5397 10489 5431 10523
rect 6101 10489 6135 10523
rect 7113 10489 7147 10523
rect 9505 10489 9539 10523
rect 12081 10489 12115 10523
rect 16589 10489 16623 10523
rect 19977 10489 20011 10523
rect 20177 10489 20211 10523
rect 21525 10489 21559 10523
rect 21741 10489 21775 10523
rect 7297 10421 7331 10455
rect 11989 10421 12023 10455
rect 12817 10421 12851 10455
rect 13277 10421 13311 10455
rect 14013 10421 14047 10455
rect 14565 10421 14599 10455
rect 17049 10421 17083 10455
rect 6377 10217 6411 10251
rect 7313 10217 7347 10251
rect 17509 10217 17543 10251
rect 17601 10217 17635 10251
rect 18245 10217 18279 10251
rect 21281 10217 21315 10251
rect 22385 10217 22419 10251
rect 3861 10149 3895 10183
rect 4077 10149 4111 10183
rect 4353 10149 4387 10183
rect 7113 10149 7147 10183
rect 8493 10149 8527 10183
rect 9197 10149 9231 10183
rect 9413 10149 9447 10183
rect 18061 10149 18095 10183
rect 22293 10149 22327 10183
rect 4997 10081 5031 10115
rect 5181 10081 5215 10115
rect 5273 10081 5307 10115
rect 5365 10081 5399 10115
rect 5549 10081 5583 10115
rect 6009 10081 6043 10115
rect 7573 10081 7607 10115
rect 7665 10081 7699 10115
rect 7849 10081 7883 10115
rect 8217 10081 8251 10115
rect 8953 10081 8987 10115
rect 11437 10081 11471 10115
rect 11989 10081 12023 10115
rect 12081 10081 12115 10115
rect 12265 10081 12299 10115
rect 12357 10081 12391 10115
rect 12541 10081 12575 10115
rect 14289 10081 14323 10115
rect 14749 10081 14783 10115
rect 14933 10081 14967 10115
rect 17233 10081 17267 10115
rect 17417 10081 17451 10115
rect 17785 10081 17819 10115
rect 17877 10081 17911 10115
rect 20729 10081 20763 10115
rect 20913 10081 20947 10115
rect 21649 10081 21683 10115
rect 22109 10081 22143 10115
rect 22753 10081 22787 10115
rect 5917 10013 5951 10047
rect 8493 10013 8527 10047
rect 8861 10013 8895 10047
rect 11529 10013 11563 10047
rect 14197 10013 14231 10047
rect 21465 10013 21499 10047
rect 21557 10013 21591 10047
rect 21741 10013 21775 10047
rect 22661 10013 22695 10047
rect 3709 9945 3743 9979
rect 4721 9945 4755 9979
rect 8309 9945 8343 9979
rect 14657 9945 14691 9979
rect 3893 9877 3927 9911
rect 4169 9877 4203 9911
rect 4353 9877 4387 9911
rect 4813 9877 4847 9911
rect 5457 9877 5491 9911
rect 7297 9877 7331 9911
rect 7481 9877 7515 9911
rect 7849 9877 7883 9911
rect 8585 9877 8619 9911
rect 8769 9877 8803 9911
rect 9045 9877 9079 9911
rect 9229 9877 9263 9911
rect 11713 9877 11747 9911
rect 12357 9877 12391 9911
rect 14749 9877 14783 9911
rect 21097 9877 21131 9911
rect 21925 9877 21959 9911
rect 22569 9877 22603 9911
rect 3341 9673 3375 9707
rect 3893 9673 3927 9707
rect 5365 9673 5399 9707
rect 5825 9673 5859 9707
rect 6101 9673 6135 9707
rect 6561 9673 6595 9707
rect 7481 9673 7515 9707
rect 14657 9673 14691 9707
rect 15485 9673 15519 9707
rect 16681 9673 16715 9707
rect 18981 9673 19015 9707
rect 19257 9673 19291 9707
rect 20729 9673 20763 9707
rect 21189 9673 21223 9707
rect 22845 9673 22879 9707
rect 5917 9605 5951 9639
rect 6377 9605 6411 9639
rect 8217 9605 8251 9639
rect 14105 9605 14139 9639
rect 15945 9605 15979 9639
rect 20821 9605 20855 9639
rect 8401 9537 8435 9571
rect 8861 9537 8895 9571
rect 9321 9537 9355 9571
rect 11437 9537 11471 9571
rect 13645 9537 13679 9571
rect 14473 9537 14507 9571
rect 14933 9537 14967 9571
rect 15577 9537 15611 9571
rect 18061 9537 18095 9571
rect 20361 9537 20395 9571
rect 3249 9469 3283 9503
rect 3433 9469 3467 9503
rect 3985 9469 4019 9503
rect 4252 9469 4286 9503
rect 5457 9469 5491 9503
rect 5641 9469 5675 9503
rect 7297 9469 7331 9503
rect 7481 9469 7515 9503
rect 7941 9469 7975 9503
rect 8033 9469 8067 9503
rect 8769 9469 8803 9503
rect 9413 9469 9447 9503
rect 11345 9469 11379 9503
rect 13737 9469 13771 9503
rect 14381 9469 14415 9503
rect 15025 9469 15059 9503
rect 15761 9469 15795 9503
rect 16129 9469 16163 9503
rect 16405 9469 16439 9503
rect 19441 9469 19475 9503
rect 20545 9469 20579 9503
rect 21465 9469 21499 9503
rect 3525 9401 3559 9435
rect 3709 9401 3743 9435
rect 6069 9401 6103 9435
rect 6285 9401 6319 9435
rect 6529 9401 6563 9435
rect 6745 9401 6779 9435
rect 8217 9401 8251 9435
rect 15485 9401 15519 9435
rect 16221 9401 16255 9435
rect 17794 9401 17828 9435
rect 19165 9401 19199 9435
rect 19625 9401 19659 9435
rect 21710 9401 21744 9435
rect 7665 9333 7699 9367
rect 9781 9333 9815 9367
rect 11713 9333 11747 9367
rect 15393 9333 15427 9367
rect 16589 9333 16623 9367
rect 18797 9333 18831 9367
rect 18965 9333 18999 9367
rect 21189 9333 21223 9367
rect 21373 9333 21407 9367
rect 5273 9129 5307 9163
rect 7205 9129 7239 9163
rect 9413 9129 9447 9163
rect 12725 9129 12759 9163
rect 16773 9129 16807 9163
rect 19901 9129 19935 9163
rect 20453 9129 20487 9163
rect 21097 9129 21131 9163
rect 22661 9129 22695 9163
rect 3884 9061 3918 9095
rect 5365 9061 5399 9095
rect 8953 9061 8987 9095
rect 12265 9061 12299 9095
rect 14749 9061 14783 9095
rect 16497 9061 16531 9095
rect 16957 9061 16991 9095
rect 17569 9061 17603 9095
rect 17785 9061 17819 9095
rect 18788 9061 18822 9095
rect 19993 9061 20027 9095
rect 20545 9061 20579 9095
rect 5457 8993 5491 9027
rect 5825 8993 5859 9027
rect 6092 8993 6126 9027
rect 8401 8993 8435 9027
rect 9229 8993 9263 9027
rect 11161 8993 11195 9027
rect 11805 8993 11839 9027
rect 12541 8993 12575 9027
rect 14657 8993 14691 9027
rect 14841 8993 14875 9027
rect 18521 8993 18555 9027
rect 20269 8993 20303 9027
rect 20729 8993 20763 9027
rect 20821 8993 20855 9027
rect 20913 8993 20947 9027
rect 21537 8993 21571 9027
rect 3617 8925 3651 8959
rect 5089 8925 5123 8959
rect 8309 8925 8343 8959
rect 9045 8925 9079 8959
rect 11069 8925 11103 8959
rect 11713 8925 11747 8959
rect 12357 8925 12391 8959
rect 16313 8925 16347 8959
rect 20177 8925 20211 8959
rect 21281 8925 21315 8959
rect 4997 8857 5031 8891
rect 8769 8857 8803 8891
rect 11529 8857 11563 8891
rect 12173 8857 12207 8891
rect 14473 8857 14507 8891
rect 17325 8857 17359 8891
rect 17417 8857 17451 8891
rect 5641 8789 5675 8823
rect 8953 8789 8987 8823
rect 12265 8789 12299 8823
rect 15025 8789 15059 8823
rect 16957 8789 16991 8823
rect 17601 8789 17635 8823
rect 20269 8789 20303 8823
rect 5917 8585 5951 8619
rect 6101 8585 6135 8619
rect 11069 8585 11103 8619
rect 13921 8585 13955 8619
rect 14565 8585 14599 8619
rect 17785 8585 17819 8619
rect 20085 8585 20119 8619
rect 20361 8585 20395 8619
rect 21373 8585 21407 8619
rect 22569 8585 22603 8619
rect 5549 8517 5583 8551
rect 6193 8517 6227 8551
rect 10885 8517 10919 8551
rect 11897 8517 11931 8551
rect 13737 8517 13771 8551
rect 14933 8517 14967 8551
rect 20729 8517 20763 8551
rect 22385 8517 22419 8551
rect 16313 8449 16347 8483
rect 16405 8449 16439 8483
rect 18705 8449 18739 8483
rect 6561 8381 6595 8415
rect 7941 8381 7975 8415
rect 8125 8381 8159 8415
rect 8217 8381 8251 8415
rect 9045 8381 9079 8415
rect 11437 8381 11471 8415
rect 11621 8381 11655 8415
rect 12081 8381 12115 8415
rect 13185 8381 13219 8415
rect 13369 8381 13403 8415
rect 14289 8381 14323 8415
rect 17877 8381 17911 8415
rect 18061 8381 18095 8415
rect 18337 8381 18371 8415
rect 20913 8381 20947 8415
rect 21097 8381 21131 8415
rect 21741 8381 21775 8415
rect 22017 8381 22051 8415
rect 22293 8381 22327 8415
rect 6377 8313 6411 8347
rect 8401 8313 8435 8347
rect 8585 8313 8619 8347
rect 11253 8313 11287 8347
rect 14381 8313 14415 8347
rect 14581 8313 14615 8347
rect 16046 8313 16080 8347
rect 16672 8313 16706 8347
rect 18521 8313 18555 8347
rect 18950 8313 18984 8347
rect 20361 8313 20395 8347
rect 21833 8313 21867 8347
rect 22201 8313 22235 8347
rect 22753 8313 22787 8347
rect 5917 8245 5951 8279
rect 7757 8245 7791 8279
rect 8769 8245 8803 8279
rect 8953 8245 8987 8279
rect 11043 8245 11077 8279
rect 11805 8245 11839 8279
rect 13185 8245 13219 8279
rect 13921 8245 13955 8279
rect 14749 8245 14783 8279
rect 17969 8245 18003 8279
rect 18153 8245 18187 8279
rect 20177 8245 20211 8279
rect 21005 8245 21039 8279
rect 21189 8245 21223 8279
rect 21373 8245 21407 8279
rect 22553 8245 22587 8279
rect 7226 8041 7260 8075
rect 7389 8041 7423 8075
rect 8493 8041 8527 8075
rect 10701 8041 10735 8075
rect 11437 8041 11471 8075
rect 11529 8041 11563 8075
rect 13093 8041 13127 8075
rect 13461 8041 13495 8075
rect 15025 8041 15059 8075
rect 18797 8041 18831 8075
rect 19533 8041 19567 8075
rect 21097 8041 21131 8075
rect 22661 8041 22695 8075
rect 4261 7973 4295 8007
rect 4721 7973 4755 8007
rect 4937 7973 4971 8007
rect 7021 7973 7055 8007
rect 7849 7973 7883 8007
rect 8309 7973 8343 8007
rect 8953 7973 8987 8007
rect 9873 7973 9907 8007
rect 10089 7973 10123 8007
rect 12265 7973 12299 8007
rect 12541 7973 12575 8007
rect 12725 7973 12759 8007
rect 14666 7973 14700 8007
rect 15209 7973 15243 8007
rect 16497 7973 16531 8007
rect 16865 7973 16899 8007
rect 17109 7973 17143 8007
rect 17325 7973 17359 8007
rect 18981 7973 19015 8007
rect 19984 7973 20018 8007
rect 22753 7973 22787 8007
rect 6745 7905 6779 7939
rect 6929 7905 6963 7939
rect 7481 7905 7515 7939
rect 8125 7905 8159 7939
rect 8401 7905 8435 7939
rect 10517 7905 10551 7939
rect 10777 7927 10811 7961
rect 10977 7903 11011 7937
rect 11161 7905 11195 7939
rect 11253 7905 11287 7939
rect 11621 7905 11655 7939
rect 13001 7905 13035 7939
rect 13277 7905 13311 7939
rect 14933 7905 14967 7939
rect 16681 7905 16715 7939
rect 19349 7905 19383 7939
rect 19441 7905 19475 7939
rect 19625 7905 19659 7939
rect 21548 7905 21582 7939
rect 22937 7905 22971 7939
rect 4629 7837 4663 7871
rect 11805 7837 11839 7871
rect 11897 7837 11931 7871
rect 19717 7837 19751 7871
rect 21281 7837 21315 7871
rect 8677 7769 8711 7803
rect 9321 7769 9355 7803
rect 13553 7769 13587 7803
rect 15577 7769 15611 7803
rect 16957 7769 16991 7803
rect 4077 7701 4111 7735
rect 4261 7701 4295 7735
rect 4905 7701 4939 7735
rect 5089 7701 5123 7735
rect 6837 7701 6871 7735
rect 7205 7701 7239 7735
rect 7849 7701 7883 7735
rect 8033 7701 8067 7735
rect 8769 7701 8803 7735
rect 8953 7701 8987 7735
rect 10057 7701 10091 7735
rect 10241 7701 10275 7735
rect 10333 7701 10367 7735
rect 11069 7701 11103 7735
rect 12265 7701 12299 7735
rect 12449 7701 12483 7735
rect 15209 7701 15243 7735
rect 17141 7701 17175 7735
rect 18981 7701 19015 7735
rect 3525 7497 3559 7531
rect 3893 7497 3927 7531
rect 5641 7497 5675 7531
rect 6561 7497 6595 7531
rect 8217 7497 8251 7531
rect 9781 7497 9815 7531
rect 11253 7497 11287 7531
rect 11345 7497 11379 7531
rect 13185 7497 13219 7531
rect 14933 7497 14967 7531
rect 15393 7497 15427 7531
rect 19257 7497 19291 7531
rect 21649 7497 21683 7531
rect 21833 7497 21867 7531
rect 6745 7429 6779 7463
rect 9873 7361 9907 7395
rect 19625 7361 19659 7395
rect 3433 7293 3467 7327
rect 3617 7293 3651 7327
rect 4169 7293 4203 7327
rect 4425 7293 4459 7327
rect 6837 7293 6871 7327
rect 8401 7293 8435 7327
rect 12458 7293 12492 7327
rect 12725 7293 12759 7327
rect 13553 7293 13587 7327
rect 15025 7293 15059 7327
rect 15209 7293 15243 7327
rect 19441 7293 19475 7327
rect 21005 7293 21039 7327
rect 21189 7293 21223 7327
rect 21281 7293 21315 7327
rect 21373 7293 21407 7327
rect 3709 7225 3743 7259
rect 3925 7225 3959 7259
rect 5825 7225 5859 7259
rect 6009 7225 6043 7259
rect 6377 7225 6411 7259
rect 7082 7225 7116 7259
rect 8668 7225 8702 7259
rect 10140 7225 10174 7259
rect 13001 7225 13035 7259
rect 13798 7225 13832 7259
rect 21925 7225 21959 7259
rect 4077 7157 4111 7191
rect 5549 7157 5583 7191
rect 6577 7157 6611 7191
rect 13201 7157 13235 7191
rect 13369 7157 13403 7191
rect 4169 6953 4203 6987
rect 5641 6953 5675 6987
rect 6193 6953 6227 6987
rect 7021 6953 7055 6987
rect 7573 6953 7607 6987
rect 10241 6953 10275 6987
rect 12357 6953 12391 6987
rect 13369 6953 13403 6987
rect 6101 6885 6135 6919
rect 7205 6885 7239 6919
rect 7389 6885 7423 6919
rect 10425 6885 10459 6919
rect 13553 6885 13587 6919
rect 3893 6817 3927 6851
rect 3985 6817 4019 6851
rect 4517 6817 4551 6851
rect 5825 6817 5859 6851
rect 6009 6817 6043 6851
rect 8686 6817 8720 6851
rect 8953 6817 8987 6851
rect 10793 6817 10827 6851
rect 10977 6817 11011 6851
rect 11233 6817 11267 6851
rect 13737 6817 13771 6851
rect 3065 6749 3099 6783
rect 3709 6749 3743 6783
rect 3801 6749 3835 6783
rect 4261 6749 4295 6783
rect 6377 6749 6411 6783
rect 3433 6681 3467 6715
rect 3525 6613 3559 6647
rect 10425 6613 10459 6647
rect 3433 6409 3467 6443
rect 3801 6409 3835 6443
rect 4353 6409 4387 6443
rect 10425 6409 10459 6443
rect 5733 6273 5767 6307
rect 3433 6205 3467 6239
rect 3709 6205 3743 6239
rect 3985 6205 4019 6239
rect 4261 6205 4295 6239
rect 5466 6205 5500 6239
rect 10609 6205 10643 6239
rect 3525 6137 3559 6171
rect 10793 6137 10827 6171
rect 4169 6069 4203 6103
rect 5273 5865 5307 5899
rect 4138 5797 4172 5831
rect 3893 5729 3927 5763
rect 22753 4097 22787 4131
rect 22937 3961 22971 3995
<< metal1 >>
rect 552 23418 23368 23440
rect 552 23366 4322 23418
rect 4374 23366 4386 23418
rect 4438 23366 4450 23418
rect 4502 23366 4514 23418
rect 4566 23366 4578 23418
rect 4630 23366 23368 23418
rect 552 23344 23368 23366
rect 7653 23307 7711 23313
rect 7653 23304 7665 23307
rect 6472 23276 7665 23304
rect 4706 23196 4712 23248
rect 4764 23236 4770 23248
rect 4764 23208 5212 23236
rect 4764 23196 4770 23208
rect 1762 23128 1768 23180
rect 1820 23128 1826 23180
rect 5184 23177 5212 23208
rect 6472 23180 6500 23276
rect 7653 23273 7665 23276
rect 7699 23273 7711 23307
rect 7653 23267 7711 23273
rect 10502 23196 10508 23248
rect 10560 23236 10566 23248
rect 11057 23239 11115 23245
rect 11057 23236 11069 23239
rect 10560 23208 11069 23236
rect 10560 23196 10566 23208
rect 11057 23205 11069 23208
rect 11103 23205 11115 23239
rect 18693 23239 18751 23245
rect 18693 23236 18705 23239
rect 11057 23199 11115 23205
rect 18156 23208 18705 23236
rect 5077 23171 5135 23177
rect 5077 23168 5089 23171
rect 1964 23140 5089 23168
rect 1964 23041 1992 23140
rect 5077 23137 5089 23140
rect 5123 23137 5135 23171
rect 5077 23131 5135 23137
rect 5169 23171 5227 23177
rect 5169 23137 5181 23171
rect 5215 23137 5227 23171
rect 5169 23131 5227 23137
rect 5092 23100 5120 23131
rect 5350 23128 5356 23180
rect 5408 23168 5414 23180
rect 5813 23171 5871 23177
rect 5813 23168 5825 23171
rect 5408 23140 5825 23168
rect 5408 23128 5414 23140
rect 5813 23137 5825 23140
rect 5859 23137 5871 23171
rect 5813 23131 5871 23137
rect 5997 23171 6055 23177
rect 5997 23137 6009 23171
rect 6043 23137 6055 23171
rect 5997 23131 6055 23137
rect 6012 23100 6040 23131
rect 6454 23128 6460 23180
rect 6512 23128 6518 23180
rect 6549 23171 6607 23177
rect 6549 23137 6561 23171
rect 6595 23137 6607 23171
rect 6549 23131 6607 23137
rect 6733 23171 6791 23177
rect 6733 23137 6745 23171
rect 6779 23168 6791 23171
rect 6914 23168 6920 23180
rect 6779 23140 6920 23168
rect 6779 23137 6791 23140
rect 6733 23131 6791 23137
rect 5092 23072 6040 23100
rect 6273 23103 6331 23109
rect 6273 23069 6285 23103
rect 6319 23100 6331 23103
rect 6564 23100 6592 23131
rect 6914 23128 6920 23140
rect 6972 23128 6978 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 8662 23128 8668 23180
rect 8720 23128 8726 23180
rect 8846 23128 8852 23180
rect 8904 23128 8910 23180
rect 13538 23128 13544 23180
rect 13596 23128 13602 23180
rect 16482 23128 16488 23180
rect 16540 23128 16546 23180
rect 7466 23100 7472 23112
rect 6319 23072 7472 23100
rect 6319 23069 6331 23072
rect 6273 23063 6331 23069
rect 7466 23060 7472 23072
rect 7524 23100 7530 23112
rect 8294 23100 8300 23112
rect 7524 23072 8300 23100
rect 7524 23060 7530 23072
rect 8294 23060 8300 23072
rect 8352 23100 8358 23112
rect 9214 23100 9220 23112
rect 8352 23072 9220 23100
rect 8352 23060 8358 23072
rect 9214 23060 9220 23072
rect 9272 23100 9278 23112
rect 9490 23100 9496 23112
rect 9272 23072 9496 23100
rect 9272 23060 9278 23072
rect 9490 23060 9496 23072
rect 9548 23060 9554 23112
rect 10134 23060 10140 23112
rect 10192 23100 10198 23112
rect 13725 23103 13783 23109
rect 13725 23100 13737 23103
rect 10192 23072 13737 23100
rect 10192 23060 10198 23072
rect 13725 23069 13737 23072
rect 13771 23100 13783 23103
rect 15286 23100 15292 23112
rect 13771 23072 15292 23100
rect 13771 23069 13783 23072
rect 13725 23063 13783 23069
rect 15286 23060 15292 23072
rect 15344 23060 15350 23112
rect 18156 23044 18184 23208
rect 18693 23205 18705 23208
rect 18739 23205 18751 23239
rect 18693 23199 18751 23205
rect 18874 23196 18880 23248
rect 18932 23245 18938 23248
rect 18932 23239 18951 23245
rect 18939 23236 18951 23239
rect 19705 23239 19763 23245
rect 19705 23236 19717 23239
rect 18939 23208 19717 23236
rect 18939 23205 18951 23208
rect 18932 23199 18951 23205
rect 19705 23205 19717 23208
rect 19751 23236 19763 23239
rect 20070 23236 20076 23248
rect 19751 23208 20076 23236
rect 19751 23205 19763 23208
rect 19705 23199 19763 23205
rect 18932 23196 18938 23199
rect 20070 23196 20076 23208
rect 20128 23196 20134 23248
rect 20254 23196 20260 23248
rect 20312 23236 20318 23248
rect 20898 23245 20904 23248
rect 20625 23239 20683 23245
rect 20625 23236 20637 23239
rect 20312 23208 20637 23236
rect 20312 23196 20318 23208
rect 20625 23205 20637 23208
rect 20671 23205 20683 23239
rect 20625 23199 20683 23205
rect 20841 23239 20904 23245
rect 20841 23205 20853 23239
rect 20887 23205 20904 23239
rect 20841 23199 20904 23205
rect 20898 23196 20904 23199
rect 20956 23196 20962 23248
rect 19058 23128 19064 23180
rect 19116 23168 19122 23180
rect 19153 23171 19211 23177
rect 19153 23168 19165 23171
rect 19116 23140 19165 23168
rect 19116 23128 19122 23140
rect 19153 23137 19165 23140
rect 19199 23137 19211 23171
rect 19153 23131 19211 23137
rect 19242 23128 19248 23180
rect 19300 23168 19306 23180
rect 19337 23171 19395 23177
rect 19337 23168 19349 23171
rect 19300 23140 19349 23168
rect 19300 23128 19306 23140
rect 19337 23137 19349 23140
rect 19383 23137 19395 23171
rect 19337 23131 19395 23137
rect 19426 23128 19432 23180
rect 19484 23128 19490 23180
rect 21174 23128 21180 23180
rect 21232 23168 21238 23180
rect 21269 23171 21327 23177
rect 21269 23168 21281 23171
rect 21232 23140 21281 23168
rect 21232 23128 21238 23140
rect 21269 23137 21281 23140
rect 21315 23137 21327 23171
rect 21269 23131 21327 23137
rect 21450 23128 21456 23180
rect 21508 23128 21514 23180
rect 22278 23128 22284 23180
rect 22336 23168 22342 23180
rect 22373 23171 22431 23177
rect 22373 23168 22385 23171
rect 22336 23140 22385 23168
rect 22336 23128 22342 23140
rect 22373 23137 22385 23140
rect 22419 23137 22431 23171
rect 22373 23131 22431 23137
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 22557 23103 22615 23109
rect 22557 23100 22569 23103
rect 20864 23072 22569 23100
rect 20864 23060 20870 23072
rect 22557 23069 22569 23072
rect 22603 23100 22615 23103
rect 22646 23100 22652 23112
rect 22603 23072 22652 23100
rect 22603 23069 22615 23072
rect 22557 23063 22615 23069
rect 22646 23060 22652 23072
rect 22704 23060 22710 23112
rect 1949 23035 2007 23041
rect 1949 23001 1961 23035
rect 1995 23001 2007 23035
rect 1949 22995 2007 23001
rect 6641 23035 6699 23041
rect 6641 23001 6653 23035
rect 6687 23032 6699 23035
rect 8110 23032 8116 23044
rect 6687 23004 8116 23032
rect 6687 23001 6699 23004
rect 6641 22995 6699 23001
rect 8110 22992 8116 23004
rect 8168 22992 8174 23044
rect 9030 22992 9036 23044
rect 9088 22992 9094 23044
rect 18138 23032 18144 23044
rect 14936 23004 18144 23032
rect 14936 22976 14964 23004
rect 18138 22992 18144 23004
rect 18196 22992 18202 23044
rect 20714 23032 20720 23044
rect 18892 23004 20720 23032
rect 4890 22924 4896 22976
rect 4948 22924 4954 22976
rect 5350 22924 5356 22976
rect 5408 22924 5414 22976
rect 11330 22924 11336 22976
rect 11388 22964 11394 22976
rect 14918 22964 14924 22976
rect 11388 22936 14924 22964
rect 11388 22924 11394 22936
rect 14918 22924 14924 22936
rect 14976 22924 14982 22976
rect 16666 22924 16672 22976
rect 16724 22924 16730 22976
rect 17954 22924 17960 22976
rect 18012 22964 18018 22976
rect 18892 22973 18920 23004
rect 20714 22992 20720 23004
rect 20772 22992 20778 23044
rect 18877 22967 18935 22973
rect 18877 22964 18889 22967
rect 18012 22936 18889 22964
rect 18012 22924 18018 22936
rect 18877 22933 18889 22936
rect 18923 22933 18935 22967
rect 18877 22927 18935 22933
rect 19058 22924 19064 22976
rect 19116 22924 19122 22976
rect 19150 22924 19156 22976
rect 19208 22924 19214 22976
rect 20162 22924 20168 22976
rect 20220 22964 20226 22976
rect 20809 22967 20867 22973
rect 20809 22964 20821 22967
rect 20220 22936 20821 22964
rect 20220 22924 20226 22936
rect 20809 22933 20821 22936
rect 20855 22933 20867 22967
rect 20809 22927 20867 22933
rect 20993 22967 21051 22973
rect 20993 22933 21005 22967
rect 21039 22964 21051 22967
rect 21174 22964 21180 22976
rect 21039 22936 21180 22964
rect 21039 22933 21051 22936
rect 20993 22927 21051 22933
rect 21174 22924 21180 22936
rect 21232 22924 21238 22976
rect 21634 22924 21640 22976
rect 21692 22924 21698 22976
rect 552 22874 23368 22896
rect 552 22822 3662 22874
rect 3714 22822 3726 22874
rect 3778 22822 3790 22874
rect 3842 22822 3854 22874
rect 3906 22822 3918 22874
rect 3970 22822 23368 22874
rect 552 22800 23368 22822
rect 6914 22760 6920 22772
rect 5276 22732 6920 22760
rect 4706 22652 4712 22704
rect 4764 22692 4770 22704
rect 4890 22692 4896 22704
rect 4764 22664 4896 22692
rect 4764 22652 4770 22664
rect 4890 22652 4896 22664
rect 4948 22652 4954 22704
rect 5276 22633 5304 22732
rect 6914 22720 6920 22732
rect 6972 22760 6978 22772
rect 8021 22763 8079 22769
rect 6972 22732 7604 22760
rect 6972 22720 6978 22732
rect 5261 22627 5319 22633
rect 5261 22593 5273 22627
rect 5307 22593 5319 22627
rect 5261 22587 5319 22593
rect 7576 22568 7604 22732
rect 8021 22729 8033 22763
rect 8067 22760 8079 22763
rect 8202 22760 8208 22772
rect 8067 22732 8208 22760
rect 8067 22729 8079 22732
rect 8021 22723 8079 22729
rect 8202 22720 8208 22732
rect 8260 22720 8266 22772
rect 8662 22720 8668 22772
rect 8720 22760 8726 22772
rect 9306 22760 9312 22772
rect 8720 22732 9312 22760
rect 8720 22720 8726 22732
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 9769 22763 9827 22769
rect 9769 22729 9781 22763
rect 9815 22760 9827 22763
rect 12158 22760 12164 22772
rect 9815 22732 12164 22760
rect 9815 22729 9827 22732
rect 9769 22723 9827 22729
rect 12158 22720 12164 22732
rect 12216 22760 12222 22772
rect 12529 22763 12587 22769
rect 12529 22760 12541 22763
rect 12216 22732 12541 22760
rect 12216 22720 12222 22732
rect 12529 22729 12541 22732
rect 12575 22729 12587 22763
rect 12529 22723 12587 22729
rect 12802 22720 12808 22772
rect 12860 22720 12866 22772
rect 15194 22720 15200 22772
rect 15252 22760 15258 22772
rect 15473 22763 15531 22769
rect 15473 22760 15485 22763
rect 15252 22732 15485 22760
rect 15252 22720 15258 22732
rect 15473 22729 15485 22732
rect 15519 22760 15531 22763
rect 15519 22732 16252 22760
rect 15519 22729 15531 22732
rect 15473 22723 15531 22729
rect 7745 22695 7803 22701
rect 7745 22661 7757 22695
rect 7791 22692 7803 22695
rect 8478 22692 8484 22704
rect 7791 22664 8484 22692
rect 7791 22661 7803 22664
rect 7745 22655 7803 22661
rect 8478 22652 8484 22664
rect 8536 22692 8542 22704
rect 8536 22664 8984 22692
rect 8536 22652 8542 22664
rect 8202 22624 8208 22636
rect 7760 22596 8208 22624
rect 4617 22559 4675 22565
rect 4617 22525 4629 22559
rect 4663 22556 4675 22559
rect 4798 22556 4804 22568
rect 4663 22528 4804 22556
rect 4663 22525 4675 22528
rect 4617 22519 4675 22525
rect 4798 22516 4804 22528
rect 4856 22516 4862 22568
rect 4893 22559 4951 22565
rect 4893 22525 4905 22559
rect 4939 22556 4951 22559
rect 5350 22556 5356 22568
rect 4939 22528 5356 22556
rect 4939 22525 4951 22528
rect 4893 22519 4951 22525
rect 4246 22448 4252 22500
rect 4304 22488 4310 22500
rect 4908 22488 4936 22519
rect 5350 22516 5356 22528
rect 5408 22516 5414 22568
rect 5902 22516 5908 22568
rect 5960 22516 5966 22568
rect 6362 22516 6368 22568
rect 6420 22516 6426 22568
rect 7466 22516 7472 22568
rect 7524 22516 7530 22568
rect 7558 22516 7564 22568
rect 7616 22516 7622 22568
rect 7760 22565 7788 22596
rect 8202 22584 8208 22596
rect 8260 22584 8266 22636
rect 7745 22559 7803 22565
rect 7745 22525 7757 22559
rect 7791 22525 7803 22559
rect 7745 22519 7803 22525
rect 7190 22488 7196 22500
rect 4304 22460 4936 22488
rect 7038 22460 7196 22488
rect 4304 22448 4310 22460
rect 7190 22448 7196 22460
rect 7248 22488 7254 22500
rect 7760 22488 7788 22519
rect 8018 22516 8024 22568
rect 8076 22556 8082 22568
rect 8481 22559 8539 22565
rect 8481 22556 8493 22559
rect 8076 22528 8493 22556
rect 8076 22516 8082 22528
rect 8481 22525 8493 22528
rect 8527 22525 8539 22559
rect 8481 22519 8539 22525
rect 8665 22559 8723 22565
rect 8665 22525 8677 22559
rect 8711 22525 8723 22559
rect 8665 22519 8723 22525
rect 7248 22460 7788 22488
rect 7837 22491 7895 22497
rect 7248 22448 7254 22460
rect 7837 22457 7849 22491
rect 7883 22457 7895 22491
rect 8294 22488 8300 22500
rect 7837 22451 7895 22457
rect 8128 22460 8300 22488
rect 7558 22380 7564 22432
rect 7616 22420 7622 22432
rect 7852 22420 7880 22451
rect 7616 22392 7880 22420
rect 8042 22423 8100 22429
rect 7616 22380 7622 22392
rect 8042 22389 8054 22423
rect 8088 22420 8100 22423
rect 8128 22420 8156 22460
rect 8294 22448 8300 22460
rect 8352 22448 8358 22500
rect 8088 22392 8156 22420
rect 8205 22423 8263 22429
rect 8088 22389 8100 22392
rect 8042 22383 8100 22389
rect 8205 22389 8217 22423
rect 8251 22420 8263 22423
rect 8570 22420 8576 22432
rect 8251 22392 8576 22420
rect 8251 22389 8263 22392
rect 8205 22383 8263 22389
rect 8570 22380 8576 22392
rect 8628 22380 8634 22432
rect 8680 22420 8708 22519
rect 8754 22516 8760 22568
rect 8812 22516 8818 22568
rect 8846 22516 8852 22568
rect 8904 22516 8910 22568
rect 8956 22556 8984 22664
rect 9030 22652 9036 22704
rect 9088 22692 9094 22704
rect 10137 22695 10195 22701
rect 10137 22692 10149 22695
rect 9088 22664 10149 22692
rect 9088 22652 9094 22664
rect 10137 22661 10149 22664
rect 10183 22661 10195 22695
rect 10137 22655 10195 22661
rect 11241 22695 11299 22701
rect 11241 22661 11253 22695
rect 11287 22692 11299 22695
rect 11974 22692 11980 22704
rect 11287 22664 11980 22692
rect 11287 22661 11299 22664
rect 11241 22655 11299 22661
rect 11974 22652 11980 22664
rect 12032 22692 12038 22704
rect 12032 22664 12434 22692
rect 12032 22652 12038 22664
rect 9125 22627 9183 22633
rect 9125 22593 9137 22627
rect 9171 22624 9183 22627
rect 10321 22627 10379 22633
rect 9171 22596 10272 22624
rect 9171 22593 9183 22596
rect 9125 22587 9183 22593
rect 9217 22559 9275 22565
rect 9217 22556 9229 22559
rect 8956 22528 9229 22556
rect 9217 22525 9229 22528
rect 9263 22525 9275 22559
rect 9217 22519 9275 22525
rect 9306 22516 9312 22568
rect 9364 22516 9370 22568
rect 9490 22516 9496 22568
rect 9548 22516 9554 22568
rect 9582 22516 9588 22568
rect 9640 22516 9646 22568
rect 10244 22556 10272 22596
rect 10321 22593 10333 22627
rect 10367 22624 10379 22627
rect 11698 22624 11704 22636
rect 10367 22596 11704 22624
rect 10367 22593 10379 22596
rect 10321 22587 10379 22593
rect 11698 22584 11704 22596
rect 11756 22584 11762 22636
rect 10505 22559 10563 22565
rect 10505 22556 10517 22559
rect 10244 22528 10517 22556
rect 10505 22525 10517 22528
rect 10551 22525 10563 22559
rect 10505 22519 10563 22525
rect 8864 22488 8892 22516
rect 8864 22460 9352 22488
rect 9324 22432 9352 22460
rect 9858 22448 9864 22500
rect 9916 22448 9922 22500
rect 10520 22488 10548 22519
rect 10594 22516 10600 22568
rect 10652 22556 10658 22568
rect 10965 22559 11023 22565
rect 10965 22556 10977 22559
rect 10652 22528 10977 22556
rect 10652 22516 10658 22528
rect 10965 22525 10977 22528
rect 11011 22525 11023 22559
rect 12406 22556 12434 22664
rect 12894 22652 12900 22704
rect 12952 22692 12958 22704
rect 13630 22692 13636 22704
rect 12952 22664 13636 22692
rect 12952 22652 12958 22664
rect 13630 22652 13636 22664
rect 13688 22652 13694 22704
rect 15562 22652 15568 22704
rect 15620 22692 15626 22704
rect 15657 22695 15715 22701
rect 15657 22692 15669 22695
rect 15620 22664 15669 22692
rect 15620 22652 15626 22664
rect 15657 22661 15669 22664
rect 15703 22661 15715 22695
rect 15657 22655 15715 22661
rect 16224 22633 16252 22732
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 17681 22763 17739 22769
rect 17681 22760 17693 22763
rect 17276 22732 17693 22760
rect 17276 22720 17282 22732
rect 17681 22729 17693 22732
rect 17727 22729 17739 22763
rect 17681 22723 17739 22729
rect 20441 22763 20499 22769
rect 20441 22729 20453 22763
rect 20487 22760 20499 22763
rect 21450 22760 21456 22772
rect 20487 22732 21456 22760
rect 20487 22729 20499 22732
rect 20441 22723 20499 22729
rect 21450 22720 21456 22732
rect 21508 22720 21514 22772
rect 21542 22720 21548 22772
rect 21600 22720 21606 22772
rect 16482 22652 16488 22704
rect 16540 22692 16546 22704
rect 18417 22695 18475 22701
rect 16540 22664 18368 22692
rect 16540 22652 16546 22664
rect 14001 22627 14059 22633
rect 14001 22624 14013 22627
rect 13464 22596 14013 22624
rect 12805 22559 12863 22565
rect 12805 22556 12817 22559
rect 12406 22528 12817 22556
rect 10965 22519 11023 22525
rect 12805 22525 12817 22528
rect 12851 22525 12863 22559
rect 12805 22519 12863 22525
rect 12897 22559 12955 22565
rect 12897 22525 12909 22559
rect 12943 22525 12955 22559
rect 13464 22556 13492 22596
rect 14001 22593 14013 22596
rect 14047 22593 14059 22627
rect 14001 22587 14059 22593
rect 16209 22627 16267 22633
rect 16209 22593 16221 22627
rect 16255 22624 16267 22627
rect 16255 22596 17172 22624
rect 16255 22593 16267 22596
rect 16209 22587 16267 22593
rect 12897 22519 12955 22525
rect 13188 22528 13492 22556
rect 11241 22491 11299 22497
rect 11241 22488 11253 22491
rect 10520 22460 11253 22488
rect 11241 22457 11253 22460
rect 11287 22457 11299 22491
rect 11241 22451 11299 22457
rect 12342 22448 12348 22500
rect 12400 22448 12406 22500
rect 12912 22488 12940 22519
rect 12728 22460 12940 22488
rect 12728 22432 12756 22460
rect 13188 22432 13216 22528
rect 13538 22516 13544 22568
rect 13596 22516 13602 22568
rect 13630 22516 13636 22568
rect 13688 22516 13694 22568
rect 14185 22559 14243 22565
rect 14185 22525 14197 22559
rect 14231 22525 14243 22559
rect 14185 22519 14243 22525
rect 13262 22448 13268 22500
rect 13320 22488 13326 22500
rect 14200 22488 14228 22519
rect 16574 22516 16580 22568
rect 16632 22556 16638 22568
rect 17037 22559 17095 22565
rect 17037 22556 17049 22559
rect 16632 22528 17049 22556
rect 16632 22516 16638 22528
rect 17037 22525 17049 22528
rect 17083 22525 17095 22559
rect 17144 22556 17172 22596
rect 17218 22584 17224 22636
rect 17276 22624 17282 22636
rect 17405 22627 17463 22633
rect 17405 22624 17417 22627
rect 17276 22596 17417 22624
rect 17276 22584 17282 22596
rect 17405 22593 17417 22596
rect 17451 22593 17463 22627
rect 17405 22587 17463 22593
rect 17954 22584 17960 22636
rect 18012 22584 18018 22636
rect 18340 22624 18368 22664
rect 18417 22661 18429 22695
rect 18463 22692 18475 22695
rect 19242 22692 19248 22704
rect 18463 22664 19248 22692
rect 18463 22661 18475 22664
rect 18417 22655 18475 22661
rect 19242 22652 19248 22664
rect 19300 22652 19306 22704
rect 20898 22692 20904 22704
rect 20456 22664 20904 22692
rect 18509 22627 18567 22633
rect 18509 22624 18521 22627
rect 18340 22596 18521 22624
rect 18509 22593 18521 22596
rect 18555 22624 18567 22627
rect 18874 22624 18880 22636
rect 18555 22596 18880 22624
rect 18555 22593 18567 22596
rect 18509 22587 18567 22593
rect 18874 22584 18880 22596
rect 18932 22584 18938 22636
rect 19150 22584 19156 22636
rect 19208 22584 19214 22636
rect 17972 22556 18000 22584
rect 17144 22528 18000 22556
rect 17037 22519 17095 22525
rect 18138 22516 18144 22568
rect 18196 22516 18202 22568
rect 18782 22516 18788 22568
rect 18840 22556 18846 22568
rect 18969 22559 19027 22565
rect 18969 22556 18981 22559
rect 18840 22528 18981 22556
rect 18840 22516 18846 22528
rect 18969 22525 18981 22528
rect 19015 22525 19027 22559
rect 18969 22519 19027 22525
rect 19794 22516 19800 22568
rect 19852 22556 19858 22568
rect 20162 22556 20168 22568
rect 19852 22528 20168 22556
rect 19852 22516 19858 22528
rect 20162 22516 20168 22528
rect 20220 22516 20226 22568
rect 20254 22516 20260 22568
rect 20312 22516 20318 22568
rect 20456 22565 20484 22664
rect 20898 22652 20904 22664
rect 20956 22692 20962 22704
rect 21085 22695 21143 22701
rect 21085 22692 21097 22695
rect 20956 22664 21097 22692
rect 20956 22652 20962 22664
rect 21085 22661 21097 22664
rect 21131 22661 21143 22695
rect 21085 22655 21143 22661
rect 21818 22652 21824 22704
rect 21876 22692 21882 22704
rect 22005 22695 22063 22701
rect 22005 22692 22017 22695
rect 21876 22664 22017 22692
rect 21876 22652 21882 22664
rect 22005 22661 22017 22664
rect 22051 22661 22063 22695
rect 22005 22655 22063 22661
rect 20806 22584 20812 22636
rect 20864 22584 20870 22636
rect 21358 22584 21364 22636
rect 21416 22624 21422 22636
rect 21545 22627 21603 22633
rect 21545 22624 21557 22627
rect 21416 22596 21557 22624
rect 21416 22584 21422 22596
rect 21545 22593 21557 22596
rect 21591 22593 21603 22627
rect 21545 22587 21603 22593
rect 21634 22584 21640 22636
rect 21692 22624 21698 22636
rect 21729 22627 21787 22633
rect 21729 22624 21741 22627
rect 21692 22596 21741 22624
rect 21692 22584 21698 22596
rect 21729 22593 21741 22596
rect 21775 22593 21787 22627
rect 21729 22587 21787 22593
rect 20441 22559 20499 22565
rect 20441 22525 20453 22559
rect 20487 22525 20499 22559
rect 20441 22519 20499 22525
rect 20714 22516 20720 22568
rect 20772 22516 20778 22568
rect 21174 22516 21180 22568
rect 21232 22516 21238 22568
rect 21266 22516 21272 22568
rect 21324 22516 21330 22568
rect 21450 22516 21456 22568
rect 21508 22516 21514 22568
rect 13320 22460 14228 22488
rect 13320 22448 13326 22460
rect 15286 22448 15292 22500
rect 15344 22448 15350 22500
rect 16666 22448 16672 22500
rect 16724 22488 16730 22500
rect 16945 22491 17003 22497
rect 16945 22488 16957 22491
rect 16724 22460 16957 22488
rect 16724 22448 16730 22460
rect 16945 22457 16957 22460
rect 16991 22457 17003 22491
rect 16945 22451 17003 22457
rect 8938 22420 8944 22432
rect 8680 22392 8944 22420
rect 8938 22380 8944 22392
rect 8996 22380 9002 22432
rect 9306 22380 9312 22432
rect 9364 22380 9370 22432
rect 10870 22380 10876 22432
rect 10928 22380 10934 22432
rect 11054 22380 11060 22432
rect 11112 22380 11118 22432
rect 12526 22380 12532 22432
rect 12584 22429 12590 22432
rect 12584 22423 12603 22429
rect 12591 22389 12603 22423
rect 12584 22383 12603 22389
rect 12584 22380 12590 22383
rect 12710 22380 12716 22432
rect 12768 22380 12774 22432
rect 13170 22380 13176 22432
rect 13228 22380 13234 22432
rect 13906 22380 13912 22432
rect 13964 22380 13970 22432
rect 14366 22380 14372 22432
rect 14424 22380 14430 22432
rect 15499 22423 15557 22429
rect 15499 22389 15511 22423
rect 15545 22420 15557 22423
rect 15930 22420 15936 22432
rect 15545 22392 15936 22420
rect 15545 22389 15557 22392
rect 15499 22383 15557 22389
rect 15930 22380 15936 22392
rect 15988 22420 15994 22432
rect 16482 22420 16488 22432
rect 15988 22392 16488 22420
rect 15988 22380 15994 22392
rect 16482 22380 16488 22392
rect 16540 22380 16546 22432
rect 16960 22420 16988 22451
rect 17126 22448 17132 22500
rect 17184 22488 17190 22500
rect 17221 22491 17279 22497
rect 17221 22488 17233 22491
rect 17184 22460 17233 22488
rect 17184 22448 17190 22460
rect 17221 22457 17233 22460
rect 17267 22457 17279 22491
rect 17221 22451 17279 22457
rect 17310 22448 17316 22500
rect 17368 22488 17374 22500
rect 17497 22491 17555 22497
rect 17497 22488 17509 22491
rect 17368 22460 17509 22488
rect 17368 22448 17374 22460
rect 17497 22457 17509 22460
rect 17543 22457 17555 22491
rect 20346 22488 20352 22500
rect 17497 22451 17555 22457
rect 17604 22460 20352 22488
rect 17604 22420 17632 22460
rect 20346 22448 20352 22460
rect 20404 22448 20410 22500
rect 21284 22488 21312 22516
rect 21284 22460 22232 22488
rect 22204 22432 22232 22460
rect 16960 22392 17632 22420
rect 17678 22380 17684 22432
rect 17736 22429 17742 22432
rect 17736 22423 17755 22429
rect 17743 22389 17755 22423
rect 17736 22383 17755 22389
rect 17736 22380 17742 22383
rect 17862 22380 17868 22432
rect 17920 22380 17926 22432
rect 20070 22380 20076 22432
rect 20128 22420 20134 22432
rect 22094 22420 22100 22432
rect 20128 22392 22100 22420
rect 20128 22380 20134 22392
rect 22094 22380 22100 22392
rect 22152 22380 22158 22432
rect 22186 22380 22192 22432
rect 22244 22380 22250 22432
rect 552 22330 23368 22352
rect 552 22278 4322 22330
rect 4374 22278 4386 22330
rect 4438 22278 4450 22330
rect 4502 22278 4514 22330
rect 4566 22278 4578 22330
rect 4630 22278 23368 22330
rect 552 22256 23368 22278
rect 4798 22176 4804 22228
rect 4856 22216 4862 22228
rect 5261 22219 5319 22225
rect 5261 22216 5273 22219
rect 4856 22188 5273 22216
rect 4856 22176 4862 22188
rect 5261 22185 5273 22188
rect 5307 22185 5319 22219
rect 5261 22179 5319 22185
rect 8938 22176 8944 22228
rect 8996 22216 9002 22228
rect 9217 22219 9275 22225
rect 9217 22216 9229 22219
rect 8996 22188 9229 22216
rect 8996 22176 9002 22188
rect 9217 22185 9229 22188
rect 9263 22216 9275 22219
rect 9582 22216 9588 22228
rect 9263 22188 9588 22216
rect 9263 22185 9275 22188
rect 9217 22179 9275 22185
rect 9582 22176 9588 22188
rect 9640 22176 9646 22228
rect 12342 22176 12348 22228
rect 12400 22216 12406 22228
rect 12529 22219 12587 22225
rect 12529 22216 12541 22219
rect 12400 22188 12541 22216
rect 12400 22176 12406 22188
rect 12529 22185 12541 22188
rect 12575 22216 12587 22219
rect 12575 22188 13860 22216
rect 12575 22185 12587 22188
rect 12529 22179 12587 22185
rect 4246 22108 4252 22160
rect 4304 22148 4310 22160
rect 4617 22151 4675 22157
rect 4617 22148 4629 22151
rect 4304 22120 4629 22148
rect 4304 22108 4310 22120
rect 4617 22117 4629 22120
rect 4663 22117 4675 22151
rect 4617 22111 4675 22117
rect 5353 22151 5411 22157
rect 5353 22117 5365 22151
rect 5399 22148 5411 22151
rect 5626 22148 5632 22160
rect 5399 22120 5632 22148
rect 5399 22117 5411 22120
rect 5353 22111 5411 22117
rect 5626 22108 5632 22120
rect 5684 22148 5690 22160
rect 6454 22148 6460 22160
rect 5684 22120 6460 22148
rect 5684 22108 5690 22120
rect 6454 22108 6460 22120
rect 6512 22108 6518 22160
rect 6730 22108 6736 22160
rect 6788 22148 6794 22160
rect 6788 22120 7236 22148
rect 6788 22108 6794 22120
rect 7208 22092 7236 22120
rect 9030 22108 9036 22160
rect 9088 22148 9094 22160
rect 12894 22148 12900 22160
rect 9088 22120 9996 22148
rect 9088 22108 9094 22120
rect 6822 22040 6828 22092
rect 6880 22040 6886 22092
rect 7190 22040 7196 22092
rect 7248 22040 7254 22092
rect 8110 22040 8116 22092
rect 8168 22040 8174 22092
rect 8941 22083 8999 22089
rect 8941 22049 8953 22083
rect 8987 22080 8999 22083
rect 9769 22083 9827 22089
rect 9769 22080 9781 22083
rect 8987 22052 9781 22080
rect 8987 22049 8999 22052
rect 8941 22043 8999 22049
rect 9769 22049 9781 22052
rect 9815 22080 9827 22083
rect 9858 22080 9864 22092
rect 9815 22052 9864 22080
rect 9815 22049 9827 22052
rect 9769 22043 9827 22049
rect 9858 22040 9864 22052
rect 9916 22040 9922 22092
rect 9968 22089 9996 22120
rect 12452 22120 12900 22148
rect 11152 22092 11204 22098
rect 9953 22083 10011 22089
rect 9953 22049 9965 22083
rect 9999 22049 10011 22083
rect 9953 22043 10011 22049
rect 10781 22083 10839 22089
rect 10781 22049 10793 22083
rect 10827 22080 10839 22083
rect 10827 22052 11152 22080
rect 10827 22049 10839 22052
rect 10781 22043 10839 22049
rect 12069 22083 12127 22089
rect 12069 22049 12081 22083
rect 12115 22080 12127 22083
rect 12452 22080 12480 22120
rect 12894 22108 12900 22120
rect 12952 22148 12958 22160
rect 13832 22148 13860 22188
rect 13906 22176 13912 22228
rect 13964 22216 13970 22228
rect 14553 22219 14611 22225
rect 14553 22216 14565 22219
rect 13964 22188 14565 22216
rect 13964 22176 13970 22188
rect 14553 22185 14565 22188
rect 14599 22185 14611 22219
rect 14553 22179 14611 22185
rect 15102 22176 15108 22228
rect 15160 22216 15166 22228
rect 15289 22219 15347 22225
rect 15289 22216 15301 22219
rect 15160 22188 15301 22216
rect 15160 22176 15166 22188
rect 15289 22185 15301 22188
rect 15335 22185 15347 22219
rect 15289 22179 15347 22185
rect 15562 22176 15568 22228
rect 15620 22216 15626 22228
rect 16114 22216 16120 22228
rect 15620 22188 16120 22216
rect 15620 22176 15626 22188
rect 16114 22176 16120 22188
rect 16172 22176 16178 22228
rect 19150 22176 19156 22228
rect 19208 22216 19214 22228
rect 20254 22216 20260 22228
rect 19208 22188 20260 22216
rect 19208 22176 19214 22188
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 21174 22176 21180 22228
rect 21232 22216 21238 22228
rect 21232 22188 22048 22216
rect 21232 22176 21238 22188
rect 12952 22120 13032 22148
rect 13832 22120 15516 22148
rect 12952 22108 12958 22120
rect 12115 22052 12480 22080
rect 12115 22049 12127 22052
rect 12069 22043 12127 22049
rect 12526 22040 12532 22092
rect 12584 22080 12590 22092
rect 13004 22089 13032 22120
rect 12621 22083 12679 22089
rect 12621 22080 12633 22083
rect 12584 22052 12633 22080
rect 12584 22040 12590 22052
rect 12621 22049 12633 22052
rect 12667 22049 12679 22083
rect 12989 22083 13047 22089
rect 12989 22080 13001 22083
rect 12967 22052 13001 22080
rect 12621 22043 12679 22049
rect 12989 22049 13001 22052
rect 13035 22049 13047 22083
rect 12989 22043 13047 22049
rect 14918 22040 14924 22092
rect 14976 22040 14982 22092
rect 11152 22034 11204 22040
rect 4982 21972 4988 22024
rect 5040 21972 5046 22024
rect 8021 22015 8079 22021
rect 8021 22012 8033 22015
rect 7116 21984 8033 22012
rect 4706 21904 4712 21956
rect 4764 21944 4770 21956
rect 5000 21944 5028 21972
rect 4764 21916 5028 21944
rect 4764 21904 4770 21916
rect 4816 21885 4844 21916
rect 6914 21904 6920 21956
rect 6972 21944 6978 21956
rect 7116 21953 7144 21984
rect 8021 21981 8033 21984
rect 8067 21981 8079 22015
rect 8021 21975 8079 21981
rect 8294 21972 8300 22024
rect 8352 22012 8358 22024
rect 8846 22012 8852 22024
rect 8352 21984 8852 22012
rect 8352 21972 8358 21984
rect 8846 21972 8852 21984
rect 8904 21972 8910 22024
rect 9033 22015 9091 22021
rect 9033 21981 9045 22015
rect 9079 21981 9091 22015
rect 9033 21975 9091 21981
rect 7101 21947 7159 21953
rect 7101 21944 7113 21947
rect 6972 21916 7113 21944
rect 6972 21904 6978 21916
rect 7101 21913 7113 21916
rect 7147 21913 7159 21947
rect 7101 21907 7159 21913
rect 7466 21904 7472 21956
rect 7524 21944 7530 21956
rect 8110 21944 8116 21956
rect 7524 21916 8116 21944
rect 7524 21904 7530 21916
rect 8110 21904 8116 21916
rect 8168 21944 8174 21956
rect 9048 21944 9076 21975
rect 9398 21972 9404 22024
rect 9456 21972 9462 22024
rect 11238 21972 11244 22024
rect 11296 21972 11302 22024
rect 12158 21972 12164 22024
rect 12216 21972 12222 22024
rect 12345 22015 12403 22021
rect 12345 21981 12357 22015
rect 12391 22012 12403 22015
rect 13265 22015 13323 22021
rect 13265 22012 13277 22015
rect 12391 21984 13277 22012
rect 12391 21981 12403 21984
rect 12345 21975 12403 21981
rect 13265 21981 13277 21984
rect 13311 22012 13323 22015
rect 13538 22012 13544 22024
rect 13311 21984 13544 22012
rect 13311 21981 13323 21984
rect 13265 21975 13323 21981
rect 13538 21972 13544 21984
rect 13596 21972 13602 22024
rect 13814 21972 13820 22024
rect 13872 22012 13878 22024
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13872 21984 14105 22012
rect 13872 21972 13878 21984
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 14185 22015 14243 22021
rect 14185 21981 14197 22015
rect 14231 22012 14243 22015
rect 14274 22012 14280 22024
rect 14231 21984 14280 22012
rect 14231 21981 14243 21984
rect 14185 21975 14243 21981
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 15013 22015 15071 22021
rect 15013 21981 15025 22015
rect 15059 22012 15071 22015
rect 15194 22012 15200 22024
rect 15059 21984 15200 22012
rect 15059 21981 15071 21984
rect 15013 21975 15071 21981
rect 15194 21972 15200 21984
rect 15252 21972 15258 22024
rect 8168 21916 9076 21944
rect 8168 21904 8174 21916
rect 11054 21904 11060 21956
rect 11112 21944 11118 21956
rect 15381 21947 15439 21953
rect 15381 21944 15393 21947
rect 11112 21916 15393 21944
rect 11112 21904 11118 21916
rect 15381 21913 15393 21916
rect 15427 21913 15439 21947
rect 15488 21944 15516 22120
rect 16482 22108 16488 22160
rect 16540 22148 16546 22160
rect 16540 22120 16896 22148
rect 16540 22108 16546 22120
rect 15746 22040 15752 22092
rect 15804 22040 15810 22092
rect 16114 22040 16120 22092
rect 16172 22040 16178 22092
rect 16206 22040 16212 22092
rect 16264 22080 16270 22092
rect 16761 22083 16819 22089
rect 16761 22080 16773 22083
rect 16264 22052 16773 22080
rect 16264 22040 16270 22052
rect 16761 22049 16773 22052
rect 16807 22049 16819 22083
rect 16761 22043 16819 22049
rect 16868 22070 16896 22120
rect 17586 22108 17592 22160
rect 17644 22148 17650 22160
rect 19334 22148 19340 22160
rect 17644 22120 19340 22148
rect 17644 22108 17650 22120
rect 19334 22108 19340 22120
rect 19392 22108 19398 22160
rect 19981 22151 20039 22157
rect 19981 22117 19993 22151
rect 20027 22148 20039 22151
rect 20346 22148 20352 22160
rect 20027 22120 20352 22148
rect 20027 22117 20039 22120
rect 19981 22111 20039 22117
rect 20346 22108 20352 22120
rect 20404 22108 20410 22160
rect 20806 22148 20812 22160
rect 20456 22120 20812 22148
rect 16868 22042 16988 22070
rect 15654 21972 15660 22024
rect 15712 21972 15718 22024
rect 16960 22012 16988 22042
rect 17034 22040 17040 22092
rect 17092 22040 17098 22092
rect 17770 22040 17776 22092
rect 17828 22080 17834 22092
rect 17865 22083 17923 22089
rect 17865 22080 17877 22083
rect 17828 22052 17877 22080
rect 17828 22040 17834 22052
rect 17865 22049 17877 22052
rect 17911 22049 17923 22083
rect 17865 22043 17923 22049
rect 18509 22083 18567 22089
rect 18509 22049 18521 22083
rect 18555 22080 18567 22083
rect 19058 22080 19064 22092
rect 18555 22052 19064 22080
rect 18555 22049 18567 22052
rect 17494 22012 17500 22024
rect 16960 21984 17500 22012
rect 17494 21972 17500 21984
rect 17552 21972 17558 22024
rect 17972 22021 18092 22046
rect 18509 22043 18567 22049
rect 19058 22040 19064 22052
rect 19116 22040 19122 22092
rect 19242 22040 19248 22092
rect 19300 22040 19306 22092
rect 19889 22083 19947 22089
rect 19889 22049 19901 22083
rect 19935 22049 19947 22083
rect 19889 22043 19947 22049
rect 17957 22018 18092 22021
rect 17957 22015 18015 22018
rect 17957 21981 17969 22015
rect 18003 21981 18015 22015
rect 17957 21975 18015 21981
rect 18064 21944 18092 22018
rect 19334 21972 19340 22024
rect 19392 22012 19398 22024
rect 19904 22012 19932 22043
rect 20162 22040 20168 22092
rect 20220 22040 20226 22092
rect 20456 22089 20484 22120
rect 20806 22108 20812 22120
rect 20864 22108 20870 22160
rect 21358 22148 21364 22160
rect 21284 22120 21364 22148
rect 20441 22083 20499 22089
rect 20441 22080 20453 22083
rect 20272 22052 20453 22080
rect 20272 22012 20300 22052
rect 20441 22049 20453 22052
rect 20487 22049 20499 22083
rect 20441 22043 20499 22049
rect 19392 21984 20300 22012
rect 20349 22015 20407 22021
rect 19392 21972 19398 21984
rect 20349 21981 20361 22015
rect 20395 22012 20407 22015
rect 21284 22012 21312 22120
rect 21358 22108 21364 22120
rect 21416 22148 21422 22160
rect 21821 22151 21879 22157
rect 21821 22148 21833 22151
rect 21416 22120 21833 22148
rect 21416 22108 21422 22120
rect 21821 22117 21833 22120
rect 21867 22117 21879 22151
rect 21821 22111 21879 22117
rect 21450 22040 21456 22092
rect 21508 22080 21514 22092
rect 21913 22083 21971 22089
rect 21913 22080 21925 22083
rect 21508 22052 21925 22080
rect 21508 22040 21514 22052
rect 21913 22049 21925 22052
rect 21959 22049 21971 22083
rect 22020 22080 22048 22188
rect 22094 22176 22100 22228
rect 22152 22216 22158 22228
rect 22152 22188 22508 22216
rect 22152 22176 22158 22188
rect 22480 22157 22508 22188
rect 22465 22151 22523 22157
rect 22465 22117 22477 22151
rect 22511 22117 22523 22151
rect 22465 22111 22523 22117
rect 22646 22108 22652 22160
rect 22704 22108 22710 22160
rect 22097 22083 22155 22089
rect 22097 22080 22109 22083
rect 22020 22052 22109 22080
rect 21913 22043 21971 22049
rect 22097 22049 22109 22052
rect 22143 22049 22155 22083
rect 22097 22043 22155 22049
rect 20395 21984 21312 22012
rect 20395 21981 20407 21984
rect 20349 21975 20407 21981
rect 21726 21972 21732 22024
rect 21784 21972 21790 22024
rect 21928 22012 21956 22043
rect 22186 22040 22192 22092
rect 22244 22040 22250 22092
rect 22370 22040 22376 22092
rect 22428 22040 22434 22092
rect 21928 21984 22232 22012
rect 19702 21944 19708 21956
rect 15488 21916 19708 21944
rect 15381 21907 15439 21913
rect 19702 21904 19708 21916
rect 19760 21904 19766 21956
rect 21453 21947 21511 21953
rect 21453 21913 21465 21947
rect 21499 21944 21511 21947
rect 21634 21944 21640 21956
rect 21499 21916 21640 21944
rect 21499 21913 21511 21916
rect 21453 21907 21511 21913
rect 21634 21904 21640 21916
rect 21692 21904 21698 21956
rect 22204 21944 22232 21984
rect 22278 21972 22284 22024
rect 22336 21972 22342 22024
rect 22373 21947 22431 21953
rect 22373 21944 22385 21947
rect 22204 21916 22385 21944
rect 22373 21913 22385 21916
rect 22419 21913 22431 21947
rect 22373 21907 22431 21913
rect 4801 21879 4859 21885
rect 4801 21845 4813 21879
rect 4847 21845 4859 21879
rect 4801 21839 4859 21845
rect 4985 21879 5043 21885
rect 4985 21845 4997 21879
rect 5031 21876 5043 21879
rect 5442 21876 5448 21888
rect 5031 21848 5448 21876
rect 5031 21845 5043 21848
rect 4985 21839 5043 21845
rect 5442 21836 5448 21848
rect 5500 21836 5506 21888
rect 8846 21836 8852 21888
rect 8904 21876 8910 21888
rect 9306 21876 9312 21888
rect 8904 21848 9312 21876
rect 8904 21836 8910 21848
rect 9306 21836 9312 21848
rect 9364 21876 9370 21888
rect 9401 21879 9459 21885
rect 9401 21876 9413 21879
rect 9364 21848 9413 21876
rect 9364 21836 9370 21848
rect 9401 21845 9413 21848
rect 9447 21845 9459 21879
rect 9401 21839 9459 21845
rect 13906 21836 13912 21888
rect 13964 21836 13970 21888
rect 14182 21836 14188 21888
rect 14240 21876 14246 21888
rect 16301 21879 16359 21885
rect 16301 21876 16313 21879
rect 14240 21848 16313 21876
rect 14240 21836 14246 21848
rect 16301 21845 16313 21848
rect 16347 21876 16359 21879
rect 17402 21876 17408 21888
rect 16347 21848 17408 21876
rect 16347 21845 16359 21848
rect 16301 21839 16359 21845
rect 17402 21836 17408 21848
rect 17460 21836 17466 21888
rect 17589 21879 17647 21885
rect 17589 21845 17601 21879
rect 17635 21876 17647 21879
rect 17678 21876 17684 21888
rect 17635 21848 17684 21876
rect 17635 21845 17647 21848
rect 17589 21839 17647 21845
rect 17678 21836 17684 21848
rect 17736 21836 17742 21888
rect 18690 21836 18696 21888
rect 18748 21836 18754 21888
rect 18782 21836 18788 21888
rect 18840 21876 18846 21888
rect 19797 21879 19855 21885
rect 19797 21876 19809 21879
rect 18840 21848 19809 21876
rect 18840 21836 18846 21848
rect 19797 21845 19809 21848
rect 19843 21876 19855 21879
rect 20530 21876 20536 21888
rect 19843 21848 20536 21876
rect 19843 21845 19855 21848
rect 19797 21839 19855 21845
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 20990 21836 20996 21888
rect 21048 21876 21054 21888
rect 21269 21879 21327 21885
rect 21269 21876 21281 21879
rect 21048 21848 21281 21876
rect 21048 21836 21054 21848
rect 21269 21845 21281 21848
rect 21315 21845 21327 21879
rect 21269 21839 21327 21845
rect 552 21786 23368 21808
rect 552 21734 3662 21786
rect 3714 21734 3726 21786
rect 3778 21734 3790 21786
rect 3842 21734 3854 21786
rect 3906 21734 3918 21786
rect 3970 21734 23368 21786
rect 552 21712 23368 21734
rect 5442 21632 5448 21684
rect 5500 21672 5506 21684
rect 5500 21644 6960 21672
rect 5500 21632 5506 21644
rect 6822 21604 6828 21616
rect 5184 21576 6828 21604
rect 5184 21454 5212 21576
rect 6822 21564 6828 21576
rect 6880 21564 6886 21616
rect 6932 21604 6960 21644
rect 7650 21632 7656 21684
rect 7708 21672 7714 21684
rect 8754 21672 8760 21684
rect 7708 21644 8760 21672
rect 7708 21632 7714 21644
rect 8754 21632 8760 21644
rect 8812 21632 8818 21684
rect 12253 21675 12311 21681
rect 12253 21641 12265 21675
rect 12299 21672 12311 21675
rect 12529 21675 12587 21681
rect 12529 21672 12541 21675
rect 12299 21644 12541 21672
rect 12299 21641 12311 21644
rect 12253 21635 12311 21641
rect 12529 21641 12541 21644
rect 12575 21672 12587 21675
rect 12802 21672 12808 21684
rect 12575 21644 12808 21672
rect 12575 21641 12587 21644
rect 12529 21635 12587 21641
rect 12802 21632 12808 21644
rect 12860 21632 12866 21684
rect 15102 21632 15108 21684
rect 15160 21672 15166 21684
rect 16669 21675 16727 21681
rect 15160 21644 16160 21672
rect 15160 21632 15166 21644
rect 6932 21576 7788 21604
rect 5261 21471 5319 21477
rect 5261 21437 5273 21471
rect 5307 21468 5319 21471
rect 6270 21468 6276 21480
rect 5307 21440 6276 21468
rect 5307 21437 5319 21440
rect 5261 21431 5319 21437
rect 6270 21428 6276 21440
rect 6328 21428 6334 21480
rect 6730 21428 6736 21480
rect 6788 21428 6794 21480
rect 6822 21428 6828 21480
rect 6880 21468 6886 21480
rect 7285 21471 7343 21477
rect 7285 21468 7297 21471
rect 6880 21440 7297 21468
rect 6880 21428 6886 21440
rect 7285 21437 7297 21440
rect 7331 21468 7343 21471
rect 7331 21440 7512 21468
rect 7331 21437 7343 21440
rect 7285 21431 7343 21437
rect 4525 21403 4583 21409
rect 4525 21369 4537 21403
rect 4571 21369 4583 21403
rect 7374 21400 7380 21412
rect 6394 21372 7380 21400
rect 4525 21363 4583 21369
rect 4540 21332 4568 21363
rect 6840 21344 6868 21372
rect 7374 21360 7380 21372
rect 7432 21360 7438 21412
rect 4706 21332 4712 21344
rect 4540 21304 4712 21332
rect 4706 21292 4712 21304
rect 4764 21292 4770 21344
rect 6822 21292 6828 21344
rect 6880 21292 6886 21344
rect 7484 21332 7512 21440
rect 7650 21428 7656 21480
rect 7708 21428 7714 21480
rect 7760 21477 7788 21576
rect 8202 21564 8208 21616
rect 8260 21604 8266 21616
rect 9125 21607 9183 21613
rect 8260 21576 9076 21604
rect 8260 21564 8266 21576
rect 9048 21536 9076 21576
rect 9125 21573 9137 21607
rect 9171 21604 9183 21607
rect 12437 21607 12495 21613
rect 9171 21576 12020 21604
rect 9171 21573 9183 21576
rect 9125 21567 9183 21573
rect 10594 21536 10600 21548
rect 7944 21508 8984 21536
rect 9048 21508 9352 21536
rect 7944 21477 7972 21508
rect 8956 21480 8984 21508
rect 7745 21471 7803 21477
rect 7745 21437 7757 21471
rect 7791 21437 7803 21471
rect 7745 21431 7803 21437
rect 7929 21471 7987 21477
rect 7929 21437 7941 21471
rect 7975 21437 7987 21471
rect 7929 21431 7987 21437
rect 7760 21400 7788 21431
rect 8018 21428 8024 21480
rect 8076 21428 8082 21480
rect 8294 21468 8300 21480
rect 8128 21440 8300 21468
rect 8128 21400 8156 21440
rect 8294 21428 8300 21440
rect 8352 21428 8358 21480
rect 8481 21471 8539 21477
rect 8481 21437 8493 21471
rect 8527 21468 8539 21471
rect 8570 21468 8576 21480
rect 8527 21440 8576 21468
rect 8527 21437 8539 21440
rect 8481 21431 8539 21437
rect 8570 21428 8576 21440
rect 8628 21428 8634 21480
rect 8662 21428 8668 21480
rect 8720 21428 8726 21480
rect 8938 21428 8944 21480
rect 8996 21428 9002 21480
rect 9214 21428 9220 21480
rect 9272 21428 9278 21480
rect 9324 21477 9352 21508
rect 9416 21508 10600 21536
rect 9309 21471 9367 21477
rect 9309 21437 9321 21471
rect 9355 21437 9367 21471
rect 9309 21431 9367 21437
rect 7760 21372 8156 21400
rect 8205 21403 8263 21409
rect 8205 21369 8217 21403
rect 8251 21400 8263 21403
rect 9416 21400 9444 21508
rect 10594 21496 10600 21508
rect 10652 21496 10658 21548
rect 10870 21496 10876 21548
rect 10928 21496 10934 21548
rect 9490 21428 9496 21480
rect 9548 21468 9554 21480
rect 9585 21471 9643 21477
rect 9585 21468 9597 21471
rect 9548 21440 9597 21468
rect 9548 21428 9554 21440
rect 9585 21437 9597 21440
rect 9631 21468 9643 21471
rect 9953 21471 10011 21477
rect 9953 21468 9965 21471
rect 9631 21440 9965 21468
rect 9631 21437 9643 21440
rect 9585 21431 9643 21437
rect 9953 21437 9965 21440
rect 9999 21437 10011 21471
rect 9953 21431 10011 21437
rect 10134 21428 10140 21480
rect 10192 21428 10198 21480
rect 10318 21428 10324 21480
rect 10376 21428 10382 21480
rect 10410 21428 10416 21480
rect 10468 21468 10474 21480
rect 10505 21471 10563 21477
rect 10505 21468 10517 21471
rect 10468 21440 10517 21468
rect 10468 21428 10474 21440
rect 10505 21437 10517 21440
rect 10551 21437 10563 21471
rect 10505 21431 10563 21437
rect 10686 21428 10692 21480
rect 10744 21428 10750 21480
rect 10965 21471 11023 21477
rect 10965 21437 10977 21471
rect 11011 21468 11023 21471
rect 11054 21468 11060 21480
rect 11011 21440 11060 21468
rect 11011 21437 11023 21440
rect 10965 21431 11023 21437
rect 11054 21428 11060 21440
rect 11112 21428 11118 21480
rect 11146 21428 11152 21480
rect 11204 21468 11210 21480
rect 11425 21471 11483 21477
rect 11425 21468 11437 21471
rect 11204 21440 11437 21468
rect 11204 21428 11210 21440
rect 11425 21437 11437 21440
rect 11471 21437 11483 21471
rect 11425 21431 11483 21437
rect 11698 21428 11704 21480
rect 11756 21428 11762 21480
rect 11992 21477 12020 21576
rect 12437 21573 12449 21607
rect 12483 21573 12495 21607
rect 12437 21567 12495 21573
rect 14936 21576 15976 21604
rect 12342 21496 12348 21548
rect 12400 21496 12406 21548
rect 12452 21536 12480 21567
rect 13173 21539 13231 21545
rect 13173 21536 13185 21539
rect 12452 21508 13185 21536
rect 13173 21505 13185 21508
rect 13219 21536 13231 21539
rect 13262 21536 13268 21548
rect 13219 21508 13268 21536
rect 13219 21505 13231 21508
rect 13173 21499 13231 21505
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 14366 21496 14372 21548
rect 14424 21496 14430 21548
rect 14936 21480 14964 21576
rect 15010 21496 15016 21548
rect 15068 21496 15074 21548
rect 15197 21539 15255 21545
rect 15197 21505 15209 21539
rect 15243 21536 15255 21539
rect 15654 21536 15660 21548
rect 15243 21508 15660 21536
rect 15243 21505 15255 21508
rect 15197 21499 15255 21505
rect 15654 21496 15660 21508
rect 15712 21536 15718 21548
rect 15749 21539 15807 21545
rect 15749 21536 15761 21539
rect 15712 21508 15761 21536
rect 15712 21496 15718 21508
rect 15749 21505 15761 21508
rect 15795 21505 15807 21539
rect 15749 21499 15807 21505
rect 11977 21471 12035 21477
rect 11977 21437 11989 21471
rect 12023 21437 12035 21471
rect 11977 21431 12035 21437
rect 12069 21471 12127 21477
rect 12069 21437 12081 21471
rect 12115 21468 12127 21471
rect 12158 21468 12164 21480
rect 12115 21440 12164 21468
rect 12115 21437 12127 21440
rect 12069 21431 12127 21437
rect 8251 21372 9444 21400
rect 9769 21403 9827 21409
rect 8251 21369 8263 21372
rect 8205 21363 8263 21369
rect 9769 21369 9781 21403
rect 9815 21400 9827 21403
rect 10597 21403 10655 21409
rect 9815 21372 10548 21400
rect 9815 21369 9827 21372
rect 9769 21363 9827 21369
rect 9401 21335 9459 21341
rect 9401 21332 9413 21335
rect 7484 21304 9413 21332
rect 9401 21301 9413 21304
rect 9447 21332 9459 21335
rect 10318 21332 10324 21344
rect 9447 21304 10324 21332
rect 9447 21301 9459 21304
rect 9401 21295 9459 21301
rect 10318 21292 10324 21304
rect 10376 21292 10382 21344
rect 10520 21332 10548 21372
rect 10597 21369 10609 21403
rect 10643 21400 10655 21403
rect 11238 21400 11244 21412
rect 10643 21372 11244 21400
rect 10643 21369 10655 21372
rect 10597 21363 10655 21369
rect 11238 21360 11244 21372
rect 11296 21400 11302 21412
rect 11517 21403 11575 21409
rect 11517 21400 11529 21403
rect 11296 21372 11529 21400
rect 11296 21360 11302 21372
rect 11517 21369 11529 21372
rect 11563 21369 11575 21403
rect 11992 21400 12020 21431
rect 12158 21428 12164 21440
rect 12216 21428 12222 21480
rect 12250 21428 12256 21480
rect 12308 21428 12314 21480
rect 12434 21468 12440 21480
rect 12406 21428 12440 21468
rect 12492 21428 12498 21480
rect 12621 21471 12679 21477
rect 12621 21437 12633 21471
rect 12667 21468 12679 21471
rect 12710 21468 12716 21480
rect 12667 21440 12716 21468
rect 12667 21437 12679 21440
rect 12621 21431 12679 21437
rect 12710 21428 12716 21440
rect 12768 21428 12774 21480
rect 13081 21471 13139 21477
rect 13081 21437 13093 21471
rect 13127 21468 13139 21471
rect 14182 21468 14188 21480
rect 13127 21440 14188 21468
rect 13127 21437 13139 21440
rect 13081 21431 13139 21437
rect 14182 21428 14188 21440
rect 14240 21428 14246 21480
rect 14918 21428 14924 21480
rect 14976 21428 14982 21480
rect 15102 21428 15108 21480
rect 15160 21428 15166 21480
rect 15841 21471 15899 21477
rect 15841 21468 15853 21471
rect 15304 21440 15853 21468
rect 12406 21400 12434 21428
rect 11992 21372 12434 21400
rect 11517 21363 11575 21369
rect 13722 21360 13728 21412
rect 13780 21400 13786 21412
rect 15120 21400 15148 21428
rect 13780 21372 15148 21400
rect 13780 21360 13786 21372
rect 11146 21332 11152 21344
rect 10520 21304 11152 21332
rect 11146 21292 11152 21304
rect 11204 21292 11210 21344
rect 11333 21335 11391 21341
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11422 21332 11428 21344
rect 11379 21304 11428 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11422 21292 11428 21304
rect 11480 21292 11486 21344
rect 11885 21335 11943 21341
rect 11885 21301 11897 21335
rect 11931 21332 11943 21335
rect 11974 21332 11980 21344
rect 11931 21304 11980 21332
rect 11931 21301 11943 21304
rect 11885 21295 11943 21301
rect 11974 21292 11980 21304
rect 12032 21292 12038 21344
rect 12713 21335 12771 21341
rect 12713 21301 12725 21335
rect 12759 21332 12771 21335
rect 13170 21332 13176 21344
rect 12759 21304 13176 21332
rect 12759 21301 12771 21304
rect 12713 21295 12771 21301
rect 13170 21292 13176 21304
rect 13228 21292 13234 21344
rect 13354 21292 13360 21344
rect 13412 21292 13418 21344
rect 13446 21292 13452 21344
rect 13504 21332 13510 21344
rect 13541 21335 13599 21341
rect 13541 21332 13553 21335
rect 13504 21304 13553 21332
rect 13504 21292 13510 21304
rect 13541 21301 13553 21304
rect 13587 21301 13599 21335
rect 13541 21295 13599 21301
rect 13630 21292 13636 21344
rect 13688 21332 13694 21344
rect 15304 21332 15332 21440
rect 15841 21437 15853 21440
rect 15887 21437 15899 21471
rect 15948 21468 15976 21576
rect 16132 21536 16160 21644
rect 16669 21641 16681 21675
rect 16715 21672 16727 21675
rect 17310 21672 17316 21684
rect 16715 21644 17316 21672
rect 16715 21641 16727 21644
rect 16669 21635 16727 21641
rect 17310 21632 17316 21644
rect 17368 21632 17374 21684
rect 17402 21632 17408 21684
rect 17460 21672 17466 21684
rect 17460 21644 17908 21672
rect 17460 21632 17466 21644
rect 16209 21607 16267 21613
rect 16209 21573 16221 21607
rect 16255 21604 16267 21607
rect 17126 21604 17132 21616
rect 16255 21576 17132 21604
rect 16255 21573 16267 21576
rect 16209 21567 16267 21573
rect 17126 21564 17132 21576
rect 17184 21564 17190 21616
rect 17494 21564 17500 21616
rect 17552 21564 17558 21616
rect 17589 21539 17647 21545
rect 16132 21508 16528 21536
rect 16500 21477 16528 21508
rect 17589 21505 17601 21539
rect 17635 21536 17647 21539
rect 17770 21536 17776 21548
rect 17635 21508 17776 21536
rect 17635 21505 17647 21508
rect 17589 21499 17647 21505
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 16301 21471 16359 21477
rect 16301 21468 16313 21471
rect 15948 21440 16313 21468
rect 15841 21431 15899 21437
rect 16301 21437 16313 21440
rect 16347 21437 16359 21471
rect 16301 21431 16359 21437
rect 16485 21471 16543 21477
rect 16485 21437 16497 21471
rect 16531 21437 16543 21471
rect 16485 21431 16543 21437
rect 15378 21360 15384 21412
rect 15436 21360 15442 21412
rect 15562 21360 15568 21412
rect 15620 21360 15626 21412
rect 15856 21400 15884 21431
rect 16666 21428 16672 21480
rect 16724 21468 16730 21480
rect 16945 21471 17003 21477
rect 16945 21468 16957 21471
rect 16724 21440 16957 21468
rect 16724 21428 16730 21440
rect 16945 21437 16957 21440
rect 16991 21437 17003 21471
rect 16945 21431 17003 21437
rect 17129 21471 17187 21477
rect 17129 21437 17141 21471
rect 17175 21468 17187 21471
rect 17218 21468 17224 21480
rect 17175 21440 17224 21468
rect 17175 21437 17187 21440
rect 17129 21431 17187 21437
rect 17218 21428 17224 21440
rect 17276 21428 17282 21480
rect 17310 21428 17316 21480
rect 17368 21428 17374 21480
rect 17497 21471 17555 21477
rect 17497 21437 17509 21471
rect 17543 21468 17555 21471
rect 17678 21468 17684 21480
rect 17543 21440 17684 21468
rect 17543 21437 17555 21440
rect 17497 21431 17555 21437
rect 17678 21428 17684 21440
rect 17736 21428 17742 21480
rect 17880 21468 17908 21644
rect 18690 21632 18696 21684
rect 18748 21672 18754 21684
rect 21726 21672 21732 21684
rect 18748 21644 21732 21672
rect 18748 21632 18754 21644
rect 21726 21632 21732 21644
rect 21784 21632 21790 21684
rect 18233 21607 18291 21613
rect 18233 21573 18245 21607
rect 18279 21604 18291 21607
rect 21453 21607 21511 21613
rect 18279 21576 20576 21604
rect 18279 21573 18291 21576
rect 18233 21567 18291 21573
rect 18046 21496 18052 21548
rect 18104 21536 18110 21548
rect 18785 21539 18843 21545
rect 18785 21536 18797 21539
rect 18104 21508 18368 21536
rect 18104 21496 18110 21508
rect 17957 21471 18015 21477
rect 17957 21468 17969 21471
rect 17880 21440 17969 21468
rect 17957 21437 17969 21440
rect 18003 21468 18015 21471
rect 18003 21440 18092 21468
rect 18003 21437 18015 21440
rect 17957 21431 18015 21437
rect 17034 21400 17040 21412
rect 15856 21372 17040 21400
rect 17034 21360 17040 21372
rect 17092 21360 17098 21412
rect 13688 21304 15332 21332
rect 13688 21292 13694 21304
rect 16758 21292 16764 21344
rect 16816 21292 16822 21344
rect 18064 21332 18092 21440
rect 18230 21360 18236 21412
rect 18288 21360 18294 21412
rect 18340 21400 18368 21508
rect 18524 21508 18797 21536
rect 18524 21477 18552 21508
rect 18785 21505 18797 21508
rect 18831 21505 18843 21539
rect 20548 21536 20576 21576
rect 21453 21573 21465 21607
rect 21499 21604 21511 21607
rect 21542 21604 21548 21616
rect 21499 21576 21548 21604
rect 21499 21573 21511 21576
rect 21453 21567 21511 21573
rect 21542 21564 21548 21576
rect 21600 21564 21606 21616
rect 18785 21499 18843 21505
rect 20364 21508 20576 21536
rect 20364 21477 20392 21508
rect 20548 21477 20576 21508
rect 21729 21539 21787 21545
rect 21729 21505 21741 21539
rect 21775 21536 21787 21539
rect 22278 21536 22284 21548
rect 21775 21508 22284 21536
rect 21775 21505 21787 21508
rect 21729 21499 21787 21505
rect 22278 21496 22284 21508
rect 22336 21496 22342 21548
rect 18509 21471 18567 21477
rect 18509 21437 18521 21471
rect 18555 21437 18567 21471
rect 18509 21431 18567 21437
rect 18693 21471 18751 21477
rect 18693 21437 18705 21471
rect 18739 21437 18751 21471
rect 18693 21431 18751 21437
rect 20348 21471 20406 21477
rect 20348 21437 20360 21471
rect 20394 21437 20406 21471
rect 20348 21431 20406 21437
rect 20441 21471 20499 21477
rect 20441 21437 20453 21471
rect 20487 21437 20499 21471
rect 20441 21431 20499 21437
rect 20533 21471 20591 21477
rect 20533 21437 20545 21471
rect 20579 21437 20591 21471
rect 20533 21431 20591 21437
rect 20626 21471 20684 21477
rect 20626 21437 20638 21471
rect 20672 21468 20684 21471
rect 20672 21440 20705 21468
rect 20672 21437 20684 21440
rect 20626 21431 20684 21437
rect 18708 21400 18736 21431
rect 18340 21372 18736 21400
rect 20456 21400 20484 21431
rect 20640 21400 20668 21431
rect 20990 21428 20996 21480
rect 21048 21428 21054 21480
rect 21177 21471 21235 21477
rect 21177 21437 21189 21471
rect 21223 21468 21235 21471
rect 21266 21468 21272 21480
rect 21223 21440 21272 21468
rect 21223 21437 21235 21440
rect 21177 21431 21235 21437
rect 21266 21428 21272 21440
rect 21324 21428 21330 21480
rect 21085 21403 21143 21409
rect 21085 21400 21097 21403
rect 20456 21372 21097 21400
rect 21085 21369 21097 21372
rect 21131 21369 21143 21403
rect 21085 21363 21143 21369
rect 18417 21335 18475 21341
rect 18417 21332 18429 21335
rect 18064 21304 18429 21332
rect 18417 21301 18429 21304
rect 18463 21301 18475 21335
rect 18417 21295 18475 21301
rect 20070 21292 20076 21344
rect 20128 21292 20134 21344
rect 20901 21335 20959 21341
rect 20901 21301 20913 21335
rect 20947 21332 20959 21335
rect 20990 21332 20996 21344
rect 20947 21304 20996 21332
rect 20947 21301 20959 21304
rect 20901 21295 20959 21301
rect 20990 21292 20996 21304
rect 21048 21292 21054 21344
rect 21266 21292 21272 21344
rect 21324 21292 21330 21344
rect 552 21242 23368 21264
rect 552 21190 4322 21242
rect 4374 21190 4386 21242
rect 4438 21190 4450 21242
rect 4502 21190 4514 21242
rect 4566 21190 4578 21242
rect 4630 21190 23368 21242
rect 552 21168 23368 21190
rect 6730 21088 6736 21140
rect 6788 21128 6794 21140
rect 6917 21131 6975 21137
rect 6917 21128 6929 21131
rect 6788 21100 6929 21128
rect 6788 21088 6794 21100
rect 6917 21097 6929 21100
rect 6963 21097 6975 21131
rect 6917 21091 6975 21097
rect 8018 21088 8024 21140
rect 8076 21128 8082 21140
rect 8205 21131 8263 21137
rect 8205 21128 8217 21131
rect 8076 21100 8217 21128
rect 8076 21088 8082 21100
rect 8205 21097 8217 21100
rect 8251 21097 8263 21131
rect 8205 21091 8263 21097
rect 8312 21100 9536 21128
rect 5902 21020 5908 21072
rect 5960 21060 5966 21072
rect 8312 21060 8340 21100
rect 9214 21060 9220 21072
rect 5960 21032 8340 21060
rect 8404 21032 9220 21060
rect 5960 21020 5966 21032
rect 4706 20952 4712 21004
rect 4764 20992 4770 21004
rect 5445 20995 5503 21001
rect 5445 20992 5457 20995
rect 4764 20964 5457 20992
rect 4764 20952 4770 20964
rect 5445 20961 5457 20964
rect 5491 20961 5503 20995
rect 5445 20955 5503 20961
rect 5626 20952 5632 21004
rect 5684 20952 5690 21004
rect 6012 21001 6040 21032
rect 5997 20995 6055 21001
rect 5997 20961 6009 20995
rect 6043 20961 6055 20995
rect 5997 20955 6055 20961
rect 6104 20964 7236 20992
rect 6104 20933 6132 20964
rect 6089 20927 6147 20933
rect 6089 20893 6101 20927
rect 6135 20893 6147 20927
rect 6089 20887 6147 20893
rect 6362 20884 6368 20936
rect 6420 20884 6426 20936
rect 7006 20884 7012 20936
rect 7064 20884 7070 20936
rect 7208 20933 7236 20964
rect 7374 20952 7380 21004
rect 7432 20952 7438 21004
rect 7469 20995 7527 21001
rect 7469 20961 7481 20995
rect 7515 20961 7527 20995
rect 7469 20955 7527 20961
rect 7653 20995 7711 21001
rect 7653 20961 7665 20995
rect 7699 20992 7711 20995
rect 8294 20992 8300 21004
rect 7699 20964 8300 20992
rect 7699 20961 7711 20964
rect 7653 20955 7711 20961
rect 7193 20927 7251 20933
rect 7193 20893 7205 20927
rect 7239 20924 7251 20927
rect 7484 20924 7512 20955
rect 8294 20952 8300 20964
rect 8352 20952 8358 21004
rect 8404 21001 8432 21032
rect 9214 21020 9220 21032
rect 9272 21060 9278 21072
rect 9508 21060 9536 21100
rect 9582 21088 9588 21140
rect 9640 21128 9646 21140
rect 9640 21100 10180 21128
rect 9640 21088 9646 21100
rect 9766 21060 9772 21072
rect 9272 21032 9444 21060
rect 9272 21020 9278 21032
rect 8389 20995 8447 21001
rect 8389 20961 8401 20995
rect 8435 20961 8447 20995
rect 8389 20955 8447 20961
rect 8570 20952 8576 21004
rect 8628 20992 8634 21004
rect 9416 21001 9444 21032
rect 9508 21032 9772 21060
rect 9508 21001 9536 21032
rect 9766 21020 9772 21032
rect 9824 21020 9830 21072
rect 9125 20995 9183 21001
rect 9125 20992 9137 20995
rect 8628 20964 9137 20992
rect 8628 20952 8634 20964
rect 9125 20961 9137 20964
rect 9171 20961 9183 20995
rect 9125 20955 9183 20961
rect 9309 20995 9367 21001
rect 9309 20961 9321 20995
rect 9355 20961 9367 20995
rect 9309 20955 9367 20961
rect 9401 20995 9459 21001
rect 9401 20961 9413 20995
rect 9447 20961 9459 20995
rect 9401 20955 9459 20961
rect 9493 20995 9551 21001
rect 9493 20961 9505 20995
rect 9539 20961 9551 20995
rect 9493 20955 9551 20961
rect 8110 20924 8116 20936
rect 7239 20896 8116 20924
rect 7239 20893 7251 20896
rect 7193 20887 7251 20893
rect 8110 20884 8116 20896
rect 8168 20924 8174 20936
rect 8481 20927 8539 20933
rect 8481 20924 8493 20927
rect 8168 20896 8493 20924
rect 8168 20884 8174 20896
rect 8481 20893 8493 20896
rect 8527 20893 8539 20927
rect 8481 20887 8539 20893
rect 8849 20927 8907 20933
rect 8849 20893 8861 20927
rect 8895 20893 8907 20927
rect 8849 20887 8907 20893
rect 6380 20856 6408 20884
rect 6730 20856 6736 20868
rect 6380 20828 6736 20856
rect 6730 20816 6736 20828
rect 6788 20856 6794 20868
rect 8754 20856 8760 20868
rect 6788 20828 8760 20856
rect 6788 20816 6794 20828
rect 8754 20816 8760 20828
rect 8812 20816 8818 20868
rect 8864 20856 8892 20887
rect 9214 20884 9220 20936
rect 9272 20924 9278 20936
rect 9324 20924 9352 20955
rect 9674 20952 9680 21004
rect 9732 20952 9738 21004
rect 10045 20995 10103 21001
rect 10045 20961 10057 20995
rect 10091 20961 10103 20995
rect 10045 20955 10103 20961
rect 10060 20924 10088 20955
rect 9272 20896 10088 20924
rect 10152 20924 10180 21100
rect 10410 21088 10416 21140
rect 10468 21088 10474 21140
rect 13630 21128 13636 21140
rect 10520 21100 13636 21128
rect 10520 21060 10548 21100
rect 13630 21088 13636 21100
rect 13688 21088 13694 21140
rect 13740 21100 14596 21128
rect 13740 21060 13768 21100
rect 10244 21032 10548 21060
rect 10612 21032 13768 21060
rect 10244 21004 10272 21032
rect 10226 20952 10232 21004
rect 10284 20952 10290 21004
rect 10321 20995 10379 21001
rect 10321 20961 10333 20995
rect 10367 20961 10379 20995
rect 10321 20955 10379 20961
rect 10336 20924 10364 20955
rect 10502 20952 10508 21004
rect 10560 20952 10566 21004
rect 10152 20896 10364 20924
rect 9272 20884 9278 20896
rect 10410 20884 10416 20936
rect 10468 20924 10474 20936
rect 10612 20924 10640 21032
rect 13820 21004 13872 21010
rect 13722 20992 13728 21004
rect 10468 20896 10640 20924
rect 12406 20964 13728 20992
rect 10468 20884 10474 20896
rect 9398 20856 9404 20868
rect 8864 20828 9404 20856
rect 9398 20816 9404 20828
rect 9456 20856 9462 20868
rect 12406 20856 12434 20964
rect 13722 20952 13728 20964
rect 13780 20952 13786 21004
rect 14568 20992 14596 21100
rect 15286 21088 15292 21140
rect 15344 21128 15350 21140
rect 15749 21131 15807 21137
rect 15749 21128 15761 21131
rect 15344 21100 15761 21128
rect 15344 21088 15350 21100
rect 15749 21097 15761 21100
rect 15795 21097 15807 21131
rect 15749 21091 15807 21097
rect 16666 21088 16672 21140
rect 16724 21088 16730 21140
rect 17862 21088 17868 21140
rect 17920 21088 17926 21140
rect 18046 21088 18052 21140
rect 18104 21088 18110 21140
rect 20885 21131 20943 21137
rect 20885 21128 20897 21131
rect 20640 21100 20897 21128
rect 15010 21020 15016 21072
rect 15068 21060 15074 21072
rect 16209 21063 16267 21069
rect 15068 21032 16160 21060
rect 15068 21020 15074 21032
rect 15194 20992 15200 21004
rect 14568 20964 15200 20992
rect 15194 20952 15200 20964
rect 15252 20992 15258 21004
rect 15657 20995 15715 21001
rect 15657 20992 15669 20995
rect 15252 20964 15669 20992
rect 15252 20952 15258 20964
rect 15657 20961 15669 20964
rect 15703 20961 15715 20995
rect 15657 20955 15715 20961
rect 15930 20952 15936 21004
rect 15988 20952 15994 21004
rect 16132 21001 16160 21032
rect 16209 21029 16221 21063
rect 16255 21060 16267 21063
rect 17681 21063 17739 21069
rect 16255 21032 16528 21060
rect 16255 21029 16267 21032
rect 16209 21023 16267 21029
rect 16500 21001 16528 21032
rect 17681 21029 17693 21063
rect 17727 21060 17739 21063
rect 17880 21060 17908 21088
rect 20640 21069 20668 21100
rect 20885 21097 20897 21100
rect 20931 21128 20943 21131
rect 21266 21128 21272 21140
rect 20931 21100 21272 21128
rect 20931 21097 20943 21100
rect 20885 21091 20943 21097
rect 21266 21088 21272 21100
rect 21324 21088 21330 21140
rect 21376 21100 21680 21128
rect 17727 21032 17908 21060
rect 20625 21063 20683 21069
rect 17727 21029 17739 21032
rect 17681 21023 17739 21029
rect 20625 21029 20637 21063
rect 20671 21029 20683 21063
rect 20990 21060 20996 21072
rect 20625 21023 20683 21029
rect 20732 21032 20996 21060
rect 16117 20995 16175 21001
rect 16117 20961 16129 20995
rect 16163 20961 16175 20995
rect 16117 20955 16175 20961
rect 16301 20995 16359 21001
rect 16301 20961 16313 20995
rect 16347 20961 16359 20995
rect 16301 20955 16359 20961
rect 16485 20995 16543 21001
rect 16485 20961 16497 20995
rect 16531 20992 16543 20995
rect 16574 20992 16580 21004
rect 16531 20964 16580 20992
rect 16531 20961 16543 20964
rect 16485 20955 16543 20961
rect 13820 20946 13872 20952
rect 13541 20927 13599 20933
rect 13541 20893 13553 20927
rect 13587 20924 13599 20927
rect 13630 20924 13636 20936
rect 13587 20896 13636 20924
rect 13587 20893 13599 20896
rect 13541 20887 13599 20893
rect 13630 20884 13636 20896
rect 13688 20884 13694 20936
rect 14274 20884 14280 20936
rect 14332 20884 14338 20936
rect 15378 20884 15384 20936
rect 15436 20924 15442 20936
rect 16316 20924 16344 20955
rect 16574 20952 16580 20964
rect 16632 20952 16638 21004
rect 16669 20995 16727 21001
rect 16669 20961 16681 20995
rect 16715 20992 16727 20995
rect 17126 20992 17132 21004
rect 16715 20964 17132 20992
rect 16715 20961 16727 20964
rect 16669 20955 16727 20961
rect 17126 20952 17132 20964
rect 17184 20952 17190 21004
rect 17494 20952 17500 21004
rect 17552 20992 17558 21004
rect 17865 20995 17923 21001
rect 17865 20992 17877 20995
rect 17552 20964 17877 20992
rect 17552 20952 17558 20964
rect 17865 20961 17877 20964
rect 17911 20992 17923 20995
rect 18230 20992 18236 21004
rect 17911 20964 18236 20992
rect 17911 20961 17923 20964
rect 17865 20955 17923 20961
rect 18230 20952 18236 20964
rect 18288 20952 18294 21004
rect 20070 20952 20076 21004
rect 20128 20952 20134 21004
rect 20257 20995 20315 21001
rect 20257 20961 20269 20995
rect 20303 20961 20315 20995
rect 20257 20955 20315 20961
rect 17310 20924 17316 20936
rect 15436 20896 15976 20924
rect 16316 20896 17316 20924
rect 15436 20884 15442 20896
rect 9456 20828 12434 20856
rect 14292 20856 14320 20884
rect 15948 20865 15976 20896
rect 17310 20884 17316 20896
rect 17368 20884 17374 20936
rect 20272 20924 20300 20955
rect 20346 20952 20352 21004
rect 20404 20952 20410 21004
rect 20441 20995 20499 21001
rect 20441 20961 20453 20995
rect 20487 20992 20499 20995
rect 20732 20992 20760 21032
rect 20990 21020 20996 21032
rect 21048 21060 21054 21072
rect 21085 21063 21143 21069
rect 21085 21060 21097 21063
rect 21048 21032 21097 21060
rect 21048 21020 21054 21032
rect 21085 21029 21097 21032
rect 21131 21060 21143 21063
rect 21376 21060 21404 21100
rect 21131 21032 21404 21060
rect 21131 21029 21143 21032
rect 21085 21023 21143 21029
rect 21542 21020 21548 21072
rect 21600 21020 21606 21072
rect 20487 20964 20760 20992
rect 21453 20995 21511 21001
rect 20487 20961 20499 20964
rect 20441 20955 20499 20961
rect 21453 20961 21465 20995
rect 21499 20992 21511 20995
rect 21560 20992 21588 21020
rect 21652 21001 21680 21100
rect 21499 20964 21588 20992
rect 21637 20995 21695 21001
rect 21499 20961 21511 20964
rect 21453 20955 21511 20961
rect 21637 20961 21649 20995
rect 21683 20961 21695 20995
rect 21637 20955 21695 20961
rect 21729 20995 21787 21001
rect 21729 20961 21741 20995
rect 21775 20992 21787 20995
rect 22278 20992 22284 21004
rect 21775 20964 22284 20992
rect 21775 20961 21787 20964
rect 21729 20955 21787 20961
rect 20456 20924 20484 20955
rect 22278 20952 22284 20964
rect 22336 20952 22342 21004
rect 20272 20896 20484 20924
rect 21545 20927 21603 20933
rect 21545 20893 21557 20927
rect 21591 20893 21603 20927
rect 21545 20887 21603 20893
rect 15933 20859 15991 20865
rect 14292 20828 15884 20856
rect 9456 20816 9462 20828
rect 5537 20791 5595 20797
rect 5537 20757 5549 20791
rect 5583 20788 5595 20791
rect 6086 20788 6092 20800
rect 5583 20760 6092 20788
rect 5583 20757 5595 20760
rect 5537 20751 5595 20757
rect 6086 20748 6092 20760
rect 6144 20748 6150 20800
rect 6362 20748 6368 20800
rect 6420 20748 6426 20800
rect 6549 20791 6607 20797
rect 6549 20757 6561 20791
rect 6595 20788 6607 20791
rect 6638 20788 6644 20800
rect 6595 20760 6644 20788
rect 6595 20757 6607 20760
rect 6549 20751 6607 20757
rect 6638 20748 6644 20760
rect 6696 20748 6702 20800
rect 7834 20748 7840 20800
rect 7892 20748 7898 20800
rect 8294 20748 8300 20800
rect 8352 20788 8358 20800
rect 8941 20791 8999 20797
rect 8941 20788 8953 20791
rect 8352 20760 8953 20788
rect 8352 20748 8358 20760
rect 8941 20757 8953 20760
rect 8987 20757 8999 20791
rect 8941 20751 8999 20757
rect 9214 20748 9220 20800
rect 9272 20788 9278 20800
rect 9582 20788 9588 20800
rect 9272 20760 9588 20788
rect 9272 20748 9278 20760
rect 9582 20748 9588 20760
rect 9640 20748 9646 20800
rect 10045 20791 10103 20797
rect 10045 20757 10057 20791
rect 10091 20788 10103 20791
rect 10686 20788 10692 20800
rect 10091 20760 10692 20788
rect 10091 20757 10103 20760
rect 10045 20751 10103 20757
rect 10686 20748 10692 20760
rect 10744 20788 10750 20800
rect 12618 20788 12624 20800
rect 10744 20760 12624 20788
rect 10744 20748 10750 20760
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 15856 20788 15884 20828
rect 15933 20825 15945 20859
rect 15979 20856 15991 20859
rect 16206 20856 16212 20868
rect 15979 20828 16212 20856
rect 15979 20825 15991 20828
rect 15933 20819 15991 20825
rect 16206 20816 16212 20828
rect 16264 20816 16270 20868
rect 20346 20816 20352 20868
rect 20404 20856 20410 20868
rect 21560 20856 21588 20887
rect 20404 20828 21588 20856
rect 20404 20816 20410 20828
rect 18690 20788 18696 20800
rect 15856 20760 18696 20788
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 19518 20748 19524 20800
rect 19576 20788 19582 20800
rect 20165 20791 20223 20797
rect 20165 20788 20177 20791
rect 19576 20760 20177 20788
rect 19576 20748 19582 20760
rect 20165 20757 20177 20760
rect 20211 20757 20223 20791
rect 20165 20751 20223 20757
rect 20622 20748 20628 20800
rect 20680 20748 20686 20800
rect 20714 20748 20720 20800
rect 20772 20748 20778 20800
rect 20916 20797 20944 20828
rect 20901 20791 20959 20797
rect 20901 20757 20913 20791
rect 20947 20757 20959 20791
rect 20901 20751 20959 20757
rect 21266 20748 21272 20800
rect 21324 20748 21330 20800
rect 552 20698 23368 20720
rect 552 20646 3662 20698
rect 3714 20646 3726 20698
rect 3778 20646 3790 20698
rect 3842 20646 3854 20698
rect 3906 20646 3918 20698
rect 3970 20646 23368 20698
rect 552 20624 23368 20646
rect 6825 20587 6883 20593
rect 6825 20553 6837 20587
rect 6871 20584 6883 20587
rect 7006 20584 7012 20596
rect 6871 20556 7012 20584
rect 6871 20553 6883 20556
rect 6825 20547 6883 20553
rect 7006 20544 7012 20556
rect 7064 20544 7070 20596
rect 20622 20544 20628 20596
rect 20680 20544 20686 20596
rect 5077 20519 5135 20525
rect 5077 20485 5089 20519
rect 5123 20516 5135 20519
rect 7650 20516 7656 20528
rect 5123 20488 7656 20516
rect 5123 20485 5135 20488
rect 5077 20479 5135 20485
rect 7650 20476 7656 20488
rect 7708 20476 7714 20528
rect 10689 20519 10747 20525
rect 10689 20485 10701 20519
rect 10735 20516 10747 20519
rect 11606 20516 11612 20528
rect 10735 20488 11612 20516
rect 10735 20485 10747 20488
rect 10689 20479 10747 20485
rect 11606 20476 11612 20488
rect 11664 20516 11670 20528
rect 11664 20488 11836 20516
rect 11664 20476 11670 20488
rect 4632 20420 5488 20448
rect 4632 20392 4660 20420
rect 4246 20340 4252 20392
rect 4304 20380 4310 20392
rect 4433 20383 4491 20389
rect 4433 20380 4445 20383
rect 4304 20352 4445 20380
rect 4304 20340 4310 20352
rect 4433 20349 4445 20352
rect 4479 20349 4491 20383
rect 4433 20343 4491 20349
rect 4614 20340 4620 20392
rect 4672 20340 4678 20392
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20349 4767 20383
rect 4709 20343 4767 20349
rect 4724 20312 4752 20343
rect 4798 20340 4804 20392
rect 4856 20340 4862 20392
rect 4893 20383 4951 20389
rect 4893 20349 4905 20383
rect 4939 20380 4951 20383
rect 5074 20380 5080 20392
rect 4939 20352 5080 20380
rect 4939 20349 4951 20352
rect 4893 20343 4951 20349
rect 5074 20340 5080 20352
rect 5132 20340 5138 20392
rect 5460 20389 5488 20420
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 11808 20457 11836 20488
rect 10229 20451 10287 20457
rect 10229 20448 10241 20451
rect 9732 20420 10241 20448
rect 9732 20408 9738 20420
rect 10229 20417 10241 20420
rect 10275 20417 10287 20451
rect 10229 20411 10287 20417
rect 11793 20451 11851 20457
rect 11793 20417 11805 20451
rect 11839 20417 11851 20451
rect 20714 20448 20720 20460
rect 11793 20411 11851 20417
rect 20548 20420 20720 20448
rect 5445 20383 5503 20389
rect 5445 20349 5457 20383
rect 5491 20349 5503 20383
rect 5445 20343 5503 20349
rect 5626 20340 5632 20392
rect 5684 20340 5690 20392
rect 5813 20383 5871 20389
rect 5813 20349 5825 20383
rect 5859 20380 5871 20383
rect 5905 20383 5963 20389
rect 5905 20380 5917 20383
rect 5859 20352 5917 20380
rect 5859 20349 5871 20352
rect 5813 20343 5871 20349
rect 5905 20349 5917 20352
rect 5951 20349 5963 20383
rect 5905 20343 5963 20349
rect 6086 20340 6092 20392
rect 6144 20340 6150 20392
rect 6730 20340 6736 20392
rect 6788 20340 6794 20392
rect 10321 20383 10379 20389
rect 10321 20349 10333 20383
rect 10367 20380 10379 20383
rect 10962 20380 10968 20392
rect 10367 20352 10968 20380
rect 10367 20349 10379 20352
rect 10321 20343 10379 20349
rect 10962 20340 10968 20352
rect 11020 20340 11026 20392
rect 11974 20340 11980 20392
rect 12032 20340 12038 20392
rect 12618 20340 12624 20392
rect 12676 20340 12682 20392
rect 12713 20383 12771 20389
rect 12713 20349 12725 20383
rect 12759 20380 12771 20383
rect 13078 20380 13084 20392
rect 12759 20352 13084 20380
rect 12759 20349 12771 20352
rect 12713 20343 12771 20349
rect 13078 20340 13084 20352
rect 13136 20340 13142 20392
rect 19058 20340 19064 20392
rect 19116 20380 19122 20392
rect 19429 20383 19487 20389
rect 19429 20380 19441 20383
rect 19116 20352 19441 20380
rect 19116 20340 19122 20352
rect 19429 20349 19441 20352
rect 19475 20349 19487 20383
rect 19429 20343 19487 20349
rect 19518 20340 19524 20392
rect 19576 20340 19582 20392
rect 20548 20389 20576 20420
rect 20714 20408 20720 20420
rect 20772 20408 20778 20460
rect 20993 20451 21051 20457
rect 20993 20417 21005 20451
rect 21039 20448 21051 20451
rect 21266 20448 21272 20460
rect 21039 20420 21272 20448
rect 21039 20417 21051 20420
rect 20993 20411 21051 20417
rect 21266 20408 21272 20420
rect 21324 20408 21330 20460
rect 20533 20383 20591 20389
rect 20533 20349 20545 20383
rect 20579 20349 20591 20383
rect 20533 20343 20591 20349
rect 20622 20340 20628 20392
rect 20680 20340 20686 20392
rect 20806 20340 20812 20392
rect 20864 20380 20870 20392
rect 21361 20383 21419 20389
rect 21361 20380 21373 20383
rect 20864 20352 21373 20380
rect 20864 20340 20870 20352
rect 21361 20349 21373 20352
rect 21407 20349 21419 20383
rect 21361 20343 21419 20349
rect 21450 20340 21456 20392
rect 21508 20340 21514 20392
rect 21637 20383 21695 20389
rect 21637 20349 21649 20383
rect 21683 20380 21695 20383
rect 22646 20380 22652 20392
rect 21683 20352 22652 20380
rect 21683 20349 21695 20352
rect 21637 20343 21695 20349
rect 22646 20340 22652 20352
rect 22704 20340 22710 20392
rect 5166 20312 5172 20324
rect 4724 20284 5172 20312
rect 5166 20272 5172 20284
rect 5224 20272 5230 20324
rect 18966 20272 18972 20324
rect 19024 20312 19030 20324
rect 19245 20315 19303 20321
rect 19245 20312 19257 20315
rect 19024 20284 19257 20312
rect 19024 20272 19030 20284
rect 19245 20281 19257 20284
rect 19291 20281 19303 20315
rect 19245 20275 19303 20281
rect 21818 20272 21824 20324
rect 21876 20272 21882 20324
rect 22462 20272 22468 20324
rect 22520 20272 22526 20324
rect 4246 20204 4252 20256
rect 4304 20204 4310 20256
rect 5994 20204 6000 20256
rect 6052 20204 6058 20256
rect 12161 20247 12219 20253
rect 12161 20213 12173 20247
rect 12207 20244 12219 20247
rect 12526 20244 12532 20256
rect 12207 20216 12532 20244
rect 12207 20213 12219 20216
rect 12161 20207 12219 20213
rect 12526 20204 12532 20216
rect 12584 20204 12590 20256
rect 12897 20247 12955 20253
rect 12897 20213 12909 20247
rect 12943 20244 12955 20247
rect 12986 20244 12992 20256
rect 12943 20216 12992 20244
rect 12943 20213 12955 20216
rect 12897 20207 12955 20213
rect 12986 20204 12992 20216
rect 13044 20204 13050 20256
rect 19521 20247 19579 20253
rect 19521 20213 19533 20247
rect 19567 20244 19579 20247
rect 19702 20244 19708 20256
rect 19567 20216 19708 20244
rect 19567 20213 19579 20216
rect 19521 20207 19579 20213
rect 19702 20204 19708 20216
rect 19760 20204 19766 20256
rect 20898 20204 20904 20256
rect 20956 20204 20962 20256
rect 21910 20204 21916 20256
rect 21968 20204 21974 20256
rect 22002 20204 22008 20256
rect 22060 20244 22066 20256
rect 22373 20247 22431 20253
rect 22373 20244 22385 20247
rect 22060 20216 22385 20244
rect 22060 20204 22066 20216
rect 22373 20213 22385 20216
rect 22419 20213 22431 20247
rect 22373 20207 22431 20213
rect 552 20154 23368 20176
rect 552 20102 4322 20154
rect 4374 20102 4386 20154
rect 4438 20102 4450 20154
rect 4502 20102 4514 20154
rect 4566 20102 4578 20154
rect 4630 20102 23368 20154
rect 552 20080 23368 20102
rect 5074 20000 5080 20052
rect 5132 20000 5138 20052
rect 15930 20040 15936 20052
rect 12268 20012 15936 20040
rect 4065 19975 4123 19981
rect 4065 19941 4077 19975
rect 4111 19972 4123 19975
rect 4154 19972 4160 19984
rect 4111 19944 4160 19972
rect 4111 19941 4123 19944
rect 4065 19935 4123 19941
rect 4154 19932 4160 19944
rect 4212 19972 4218 19984
rect 4617 19975 4675 19981
rect 4617 19972 4629 19975
rect 4212 19944 4629 19972
rect 4212 19932 4218 19944
rect 4617 19941 4629 19944
rect 4663 19972 4675 19975
rect 4890 19972 4896 19984
rect 4663 19944 4896 19972
rect 4663 19941 4675 19944
rect 4617 19935 4675 19941
rect 4890 19932 4896 19944
rect 4948 19932 4954 19984
rect 5092 19972 5120 20000
rect 10962 19972 10968 19984
rect 5092 19944 5304 19972
rect 5166 19904 5172 19916
rect 4540 19876 5172 19904
rect 4540 19845 4568 19876
rect 5166 19864 5172 19876
rect 5224 19864 5230 19916
rect 5276 19913 5304 19944
rect 10704 19944 10968 19972
rect 5261 19907 5319 19913
rect 5261 19873 5273 19907
rect 5307 19873 5319 19907
rect 5261 19867 5319 19873
rect 5994 19864 6000 19916
rect 6052 19864 6058 19916
rect 7006 19864 7012 19916
rect 7064 19864 7070 19916
rect 10321 19907 10379 19913
rect 10321 19873 10333 19907
rect 10367 19904 10379 19907
rect 10502 19904 10508 19916
rect 10367 19876 10508 19904
rect 10367 19873 10379 19876
rect 10321 19867 10379 19873
rect 10502 19864 10508 19876
rect 10560 19864 10566 19916
rect 10704 19913 10732 19944
rect 10962 19932 10968 19944
rect 11020 19972 11026 19984
rect 11020 19944 11362 19972
rect 11020 19932 11026 19944
rect 12268 19916 12296 20012
rect 15930 20000 15936 20012
rect 15988 20000 15994 20052
rect 17954 20040 17960 20052
rect 17604 20012 17960 20040
rect 12342 19932 12348 19984
rect 12400 19972 12406 19984
rect 14550 19972 14556 19984
rect 12400 19944 14556 19972
rect 12400 19932 12406 19944
rect 14550 19932 14556 19944
rect 14608 19932 14614 19984
rect 17604 19981 17632 20012
rect 17954 20000 17960 20012
rect 18012 20040 18018 20052
rect 18230 20040 18236 20052
rect 18012 20012 18236 20040
rect 18012 20000 18018 20012
rect 18230 20000 18236 20012
rect 18288 20000 18294 20052
rect 21450 20000 21456 20052
rect 21508 20000 21514 20052
rect 17313 19975 17371 19981
rect 16408 19944 16988 19972
rect 10689 19907 10747 19913
rect 10689 19873 10701 19907
rect 10735 19873 10747 19907
rect 10689 19867 10747 19873
rect 11146 19864 11152 19916
rect 11204 19904 11210 19916
rect 11977 19907 12035 19913
rect 11977 19904 11989 19907
rect 11204 19876 11989 19904
rect 11204 19864 11210 19876
rect 11977 19873 11989 19876
rect 12023 19904 12035 19907
rect 12066 19904 12072 19916
rect 12023 19876 12072 19904
rect 12023 19873 12035 19876
rect 11977 19867 12035 19873
rect 12066 19864 12072 19876
rect 12124 19864 12130 19916
rect 12250 19864 12256 19916
rect 12308 19904 12314 19916
rect 12437 19907 12495 19913
rect 12437 19904 12449 19907
rect 12308 19876 12449 19904
rect 12308 19864 12314 19876
rect 12437 19873 12449 19876
rect 12483 19873 12495 19907
rect 12437 19867 12495 19873
rect 12618 19864 12624 19916
rect 12676 19904 12682 19916
rect 13173 19907 13231 19913
rect 13173 19904 13185 19907
rect 12676 19876 13185 19904
rect 12676 19864 12682 19876
rect 13173 19873 13185 19876
rect 13219 19873 13231 19907
rect 13633 19907 13691 19913
rect 13633 19904 13645 19907
rect 13173 19867 13231 19873
rect 13556 19876 13645 19904
rect 4525 19839 4583 19845
rect 4525 19805 4537 19839
rect 4571 19805 4583 19839
rect 4525 19799 4583 19805
rect 6086 19796 6092 19848
rect 6144 19796 6150 19848
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 7558 19836 7564 19848
rect 6779 19808 7564 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 7558 19796 7564 19808
rect 7616 19836 7622 19848
rect 8849 19839 8907 19845
rect 8849 19836 8861 19839
rect 7616 19808 8861 19836
rect 7616 19796 7622 19808
rect 8849 19805 8861 19808
rect 8895 19805 8907 19839
rect 8849 19799 8907 19805
rect 13078 19796 13084 19848
rect 13136 19796 13142 19848
rect 13556 19780 13584 19876
rect 13633 19873 13645 19876
rect 13679 19873 13691 19907
rect 13633 19867 13691 19873
rect 13771 19907 13829 19913
rect 13771 19873 13783 19907
rect 13817 19904 13829 19907
rect 13906 19904 13912 19916
rect 13817 19876 13912 19904
rect 13817 19873 13829 19876
rect 13771 19867 13829 19873
rect 13906 19864 13912 19876
rect 13964 19864 13970 19916
rect 16408 19845 16436 19944
rect 16485 19907 16543 19913
rect 16485 19873 16497 19907
rect 16531 19904 16543 19907
rect 16758 19904 16764 19916
rect 16531 19876 16764 19904
rect 16531 19873 16543 19876
rect 16485 19867 16543 19873
rect 16758 19864 16764 19876
rect 16816 19864 16822 19916
rect 16960 19913 16988 19944
rect 17313 19941 17325 19975
rect 17359 19972 17371 19975
rect 17589 19975 17647 19981
rect 17589 19972 17601 19975
rect 17359 19944 17601 19972
rect 17359 19941 17371 19944
rect 17313 19935 17371 19941
rect 17589 19941 17601 19944
rect 17635 19941 17647 19975
rect 17589 19935 17647 19941
rect 17770 19932 17776 19984
rect 17828 19981 17834 19984
rect 17828 19975 17847 19981
rect 17835 19972 17847 19975
rect 18138 19972 18144 19984
rect 17835 19944 18144 19972
rect 17835 19941 17847 19944
rect 17828 19935 17847 19941
rect 17828 19932 17834 19935
rect 18138 19932 18144 19944
rect 18196 19972 18202 19984
rect 18196 19944 18460 19972
rect 18196 19932 18202 19944
rect 18432 19913 18460 19944
rect 18506 19932 18512 19984
rect 18564 19972 18570 19984
rect 19058 19972 19064 19984
rect 18564 19944 19064 19972
rect 18564 19932 18570 19944
rect 19058 19932 19064 19944
rect 19116 19932 19122 19984
rect 20346 19972 20352 19984
rect 19812 19944 20352 19972
rect 16945 19907 17003 19913
rect 16945 19873 16957 19907
rect 16991 19873 17003 19907
rect 16945 19867 17003 19873
rect 17038 19907 17096 19913
rect 17038 19873 17050 19907
rect 17084 19873 17096 19907
rect 18325 19907 18383 19913
rect 18325 19904 18337 19907
rect 17038 19867 17096 19873
rect 17880 19876 18337 19904
rect 16393 19839 16451 19845
rect 16393 19836 16405 19839
rect 13740 19808 16405 19836
rect 4338 19728 4344 19780
rect 4396 19728 4402 19780
rect 4893 19771 4951 19777
rect 4893 19768 4905 19771
rect 4724 19740 4905 19768
rect 4246 19660 4252 19712
rect 4304 19700 4310 19712
rect 4724 19700 4752 19740
rect 4893 19737 4905 19740
rect 4939 19737 4951 19771
rect 4893 19731 4951 19737
rect 6365 19771 6423 19777
rect 6365 19737 6377 19771
rect 6411 19768 6423 19771
rect 6825 19771 6883 19777
rect 6825 19768 6837 19771
rect 6411 19740 6837 19768
rect 6411 19737 6423 19740
rect 6365 19731 6423 19737
rect 6825 19737 6837 19740
rect 6871 19768 6883 19771
rect 7098 19768 7104 19780
rect 6871 19740 7104 19768
rect 6871 19737 6883 19740
rect 6825 19731 6883 19737
rect 7098 19728 7104 19740
rect 7156 19728 7162 19780
rect 7193 19771 7251 19777
rect 7193 19737 7205 19771
rect 7239 19768 7251 19771
rect 7239 19740 12434 19768
rect 7239 19737 7251 19740
rect 7193 19731 7251 19737
rect 4304 19672 4752 19700
rect 4304 19660 4310 19672
rect 4798 19660 4804 19712
rect 4856 19700 4862 19712
rect 5169 19703 5227 19709
rect 5169 19700 5181 19703
rect 4856 19672 5181 19700
rect 4856 19660 4862 19672
rect 5169 19669 5181 19672
rect 5215 19669 5227 19703
rect 5169 19663 5227 19669
rect 5534 19660 5540 19712
rect 5592 19660 5598 19712
rect 12406 19700 12434 19740
rect 13538 19728 13544 19780
rect 13596 19728 13602 19780
rect 13740 19700 13768 19808
rect 16393 19805 16405 19808
rect 16439 19805 16451 19839
rect 16776 19836 16804 19864
rect 17052 19836 17080 19867
rect 16776 19808 17080 19836
rect 16393 19799 16451 19805
rect 16850 19728 16856 19780
rect 16908 19728 16914 19780
rect 17880 19712 17908 19876
rect 18325 19873 18337 19876
rect 18371 19873 18383 19907
rect 18325 19867 18383 19873
rect 18417 19907 18475 19913
rect 18417 19873 18429 19907
rect 18463 19873 18475 19907
rect 18966 19904 18972 19916
rect 18417 19867 18475 19873
rect 18616 19876 18972 19904
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19805 18199 19839
rect 18141 19799 18199 19805
rect 18156 19768 18184 19799
rect 18230 19796 18236 19848
rect 18288 19796 18294 19848
rect 18616 19845 18644 19876
rect 18966 19864 18972 19876
rect 19024 19864 19030 19916
rect 19245 19907 19303 19913
rect 19245 19873 19257 19907
rect 19291 19904 19303 19907
rect 19518 19904 19524 19916
rect 19291 19876 19524 19904
rect 19291 19873 19303 19876
rect 19245 19867 19303 19873
rect 19518 19864 19524 19876
rect 19576 19864 19582 19916
rect 19702 19864 19708 19916
rect 19760 19864 19766 19916
rect 19812 19845 19840 19944
rect 20346 19932 20352 19944
rect 20404 19932 20410 19984
rect 21174 19932 21180 19984
rect 21232 19972 21238 19984
rect 22002 19972 22008 19984
rect 21232 19944 22008 19972
rect 21232 19932 21238 19944
rect 22002 19932 22008 19944
rect 22060 19972 22066 19984
rect 22060 19944 22324 19972
rect 22060 19932 22066 19944
rect 20162 19864 20168 19916
rect 20220 19864 20226 19916
rect 20530 19864 20536 19916
rect 20588 19864 20594 19916
rect 20714 19864 20720 19916
rect 20772 19904 20778 19916
rect 22296 19913 22324 19944
rect 20809 19907 20867 19913
rect 20809 19904 20821 19907
rect 20772 19876 20821 19904
rect 20772 19864 20778 19876
rect 20809 19873 20821 19876
rect 20855 19873 20867 19907
rect 20809 19867 20867 19873
rect 20993 19907 21051 19913
rect 20993 19873 21005 19907
rect 21039 19904 21051 19907
rect 21450 19907 21508 19913
rect 21450 19904 21462 19907
rect 21039 19876 21462 19904
rect 21039 19873 21051 19876
rect 20993 19867 21051 19873
rect 21450 19873 21462 19876
rect 21496 19904 21508 19907
rect 22281 19907 22339 19913
rect 21496 19876 22094 19904
rect 21496 19873 21508 19876
rect 21450 19867 21508 19873
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 19429 19839 19487 19845
rect 19429 19805 19441 19839
rect 19475 19836 19487 19839
rect 19797 19839 19855 19845
rect 19797 19836 19809 19839
rect 19475 19808 19809 19836
rect 19475 19805 19487 19808
rect 19429 19799 19487 19805
rect 19797 19805 19809 19808
rect 19843 19805 19855 19839
rect 19797 19799 19855 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 18690 19768 18696 19780
rect 18156 19740 18696 19768
rect 18690 19728 18696 19740
rect 18748 19728 18754 19780
rect 19904 19768 19932 19799
rect 19978 19796 19984 19848
rect 20036 19796 20042 19848
rect 20180 19836 20208 19864
rect 20625 19839 20683 19845
rect 20180 19808 20576 19836
rect 20548 19768 20576 19808
rect 20625 19805 20637 19839
rect 20671 19836 20683 19839
rect 21266 19836 21272 19848
rect 20671 19808 21272 19836
rect 20671 19805 20683 19808
rect 20625 19799 20683 19805
rect 21266 19796 21272 19808
rect 21324 19796 21330 19848
rect 21910 19796 21916 19848
rect 21968 19796 21974 19848
rect 22066 19836 22094 19876
rect 22281 19873 22293 19907
rect 22327 19873 22339 19907
rect 22281 19867 22339 19873
rect 22370 19864 22376 19916
rect 22428 19864 22434 19916
rect 22557 19907 22615 19913
rect 22557 19873 22569 19907
rect 22603 19904 22615 19907
rect 22738 19904 22744 19916
rect 22603 19876 22744 19904
rect 22603 19873 22615 19876
rect 22557 19867 22615 19873
rect 22738 19864 22744 19876
rect 22796 19864 22802 19916
rect 22830 19836 22836 19848
rect 22066 19808 22836 19836
rect 22830 19796 22836 19808
rect 22888 19796 22894 19848
rect 23014 19796 23020 19848
rect 23072 19796 23078 19848
rect 21928 19768 21956 19796
rect 19904 19740 20392 19768
rect 20548 19740 21956 19768
rect 12406 19672 13768 19700
rect 13814 19660 13820 19712
rect 13872 19660 13878 19712
rect 17773 19703 17831 19709
rect 17773 19669 17785 19703
rect 17819 19700 17831 19703
rect 17862 19700 17868 19712
rect 17819 19672 17868 19700
rect 17819 19669 17831 19672
rect 17773 19663 17831 19669
rect 17862 19660 17868 19672
rect 17920 19660 17926 19712
rect 17957 19703 18015 19709
rect 17957 19669 17969 19703
rect 18003 19700 18015 19703
rect 18230 19700 18236 19712
rect 18003 19672 18236 19700
rect 18003 19669 18015 19672
rect 17957 19663 18015 19669
rect 18230 19660 18236 19672
rect 18288 19660 18294 19712
rect 19518 19660 19524 19712
rect 19576 19660 19582 19712
rect 20364 19709 20392 19740
rect 20349 19703 20407 19709
rect 20349 19669 20361 19703
rect 20395 19700 20407 19703
rect 20714 19700 20720 19712
rect 20395 19672 20720 19700
rect 20395 19669 20407 19672
rect 20349 19663 20407 19669
rect 20714 19660 20720 19672
rect 20772 19660 20778 19712
rect 21082 19660 21088 19712
rect 21140 19700 21146 19712
rect 21269 19703 21327 19709
rect 21269 19700 21281 19703
rect 21140 19672 21281 19700
rect 21140 19660 21146 19672
rect 21269 19669 21281 19672
rect 21315 19669 21327 19703
rect 21269 19663 21327 19669
rect 21821 19703 21879 19709
rect 21821 19669 21833 19703
rect 21867 19700 21879 19703
rect 22186 19700 22192 19712
rect 21867 19672 22192 19700
rect 21867 19669 21879 19672
rect 21821 19663 21879 19669
rect 22186 19660 22192 19672
rect 22244 19660 22250 19712
rect 552 19610 23368 19632
rect 552 19558 3662 19610
rect 3714 19558 3726 19610
rect 3778 19558 3790 19610
rect 3842 19558 3854 19610
rect 3906 19558 3918 19610
rect 3970 19558 23368 19610
rect 552 19536 23368 19558
rect 4525 19499 4583 19505
rect 4525 19465 4537 19499
rect 4571 19496 4583 19499
rect 4798 19496 4804 19508
rect 4571 19468 4804 19496
rect 4571 19465 4583 19468
rect 4525 19459 4583 19465
rect 4798 19456 4804 19468
rect 4856 19456 4862 19508
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 5261 19499 5319 19505
rect 5261 19496 5273 19499
rect 5224 19468 5273 19496
rect 5224 19456 5230 19468
rect 5261 19465 5273 19468
rect 5307 19465 5319 19499
rect 5261 19459 5319 19465
rect 9677 19499 9735 19505
rect 9677 19465 9689 19499
rect 9723 19496 9735 19499
rect 9858 19496 9864 19508
rect 9723 19468 9864 19496
rect 9723 19465 9735 19468
rect 9677 19459 9735 19465
rect 9858 19456 9864 19468
rect 9916 19456 9922 19508
rect 11977 19499 12035 19505
rect 11977 19465 11989 19499
rect 12023 19496 12035 19499
rect 13078 19496 13084 19508
rect 12023 19468 13084 19496
rect 12023 19465 12035 19468
rect 11977 19459 12035 19465
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 13357 19499 13415 19505
rect 13357 19465 13369 19499
rect 13403 19496 13415 19499
rect 14369 19499 14427 19505
rect 14369 19496 14381 19499
rect 13403 19468 14381 19496
rect 13403 19465 13415 19468
rect 13357 19459 13415 19465
rect 14369 19465 14381 19468
rect 14415 19496 14427 19499
rect 14734 19496 14740 19508
rect 14415 19468 14740 19496
rect 14415 19465 14427 19468
rect 14369 19459 14427 19465
rect 14734 19456 14740 19468
rect 14792 19456 14798 19508
rect 18690 19456 18696 19508
rect 18748 19456 18754 19508
rect 22186 19456 22192 19508
rect 22244 19456 22250 19508
rect 4816 19428 4844 19456
rect 7561 19431 7619 19437
rect 4816 19400 5396 19428
rect 4154 19320 4160 19372
rect 4212 19320 4218 19372
rect 4706 19320 4712 19372
rect 4764 19320 4770 19372
rect 5166 19320 5172 19372
rect 5224 19320 5230 19372
rect 5368 19369 5396 19400
rect 7561 19397 7573 19431
rect 7607 19428 7619 19431
rect 7607 19400 12103 19428
rect 7607 19397 7619 19400
rect 7561 19391 7619 19397
rect 5353 19363 5411 19369
rect 5353 19329 5365 19363
rect 5399 19329 5411 19363
rect 5353 19323 5411 19329
rect 7098 19320 7104 19372
rect 7156 19320 7162 19372
rect 11701 19363 11759 19369
rect 7944 19332 8156 19360
rect 4246 19252 4252 19304
rect 4304 19252 4310 19304
rect 4338 19252 4344 19304
rect 4396 19252 4402 19304
rect 4798 19252 4804 19304
rect 4856 19252 4862 19304
rect 5261 19295 5319 19301
rect 5261 19261 5273 19295
rect 5307 19292 5319 19295
rect 5442 19292 5448 19304
rect 5307 19264 5448 19292
rect 5307 19261 5319 19264
rect 5261 19255 5319 19261
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 5994 19252 6000 19304
rect 6052 19292 6058 19304
rect 6273 19295 6331 19301
rect 6273 19292 6285 19295
rect 6052 19264 6285 19292
rect 6052 19252 6058 19264
rect 6273 19261 6285 19264
rect 6319 19261 6331 19295
rect 6273 19255 6331 19261
rect 6457 19295 6515 19301
rect 6457 19261 6469 19295
rect 6503 19292 6515 19295
rect 7006 19292 7012 19304
rect 6503 19264 7012 19292
rect 6503 19261 6515 19264
rect 6457 19255 6515 19261
rect 7006 19252 7012 19264
rect 7064 19252 7070 19304
rect 7190 19252 7196 19304
rect 7248 19252 7254 19304
rect 7466 19252 7472 19304
rect 7524 19292 7530 19304
rect 7653 19295 7711 19301
rect 7653 19292 7665 19295
rect 7524 19264 7665 19292
rect 7524 19252 7530 19264
rect 7653 19261 7665 19264
rect 7699 19261 7711 19295
rect 7653 19255 7711 19261
rect 7834 19252 7840 19304
rect 7892 19292 7898 19304
rect 7944 19292 7972 19332
rect 7892 19264 7972 19292
rect 7892 19252 7898 19264
rect 8018 19252 8024 19304
rect 8076 19252 8082 19304
rect 8128 19292 8156 19332
rect 11701 19329 11713 19363
rect 11747 19360 11759 19363
rect 11974 19360 11980 19372
rect 11747 19332 11980 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 11974 19320 11980 19332
rect 12032 19320 12038 19372
rect 12075 19360 12103 19400
rect 12158 19388 12164 19440
rect 12216 19388 12222 19440
rect 12713 19431 12771 19437
rect 12713 19397 12725 19431
rect 12759 19428 12771 19431
rect 12986 19428 12992 19440
rect 12759 19400 12992 19428
rect 12759 19397 12771 19400
rect 12713 19391 12771 19397
rect 12986 19388 12992 19400
rect 13044 19388 13050 19440
rect 14921 19431 14979 19437
rect 14921 19397 14933 19431
rect 14967 19428 14979 19431
rect 18141 19431 18199 19437
rect 14967 19400 15056 19428
rect 14967 19397 14979 19400
rect 14921 19391 14979 19397
rect 12342 19360 12348 19372
rect 12075 19332 12348 19360
rect 12342 19320 12348 19332
rect 12400 19320 12406 19372
rect 12526 19320 12532 19372
rect 12584 19360 12590 19372
rect 12897 19363 12955 19369
rect 12897 19360 12909 19363
rect 12584 19332 12909 19360
rect 12584 19320 12590 19332
rect 12897 19329 12909 19332
rect 12943 19360 12955 19363
rect 13078 19360 13084 19372
rect 12943 19332 13084 19360
rect 12943 19329 12955 19332
rect 12897 19323 12955 19329
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 13633 19363 13691 19369
rect 13633 19329 13645 19363
rect 13679 19360 13691 19363
rect 13906 19360 13912 19372
rect 13679 19332 13912 19360
rect 13679 19329 13691 19332
rect 13633 19323 13691 19329
rect 13906 19320 13912 19332
rect 13964 19320 13970 19372
rect 13998 19320 14004 19372
rect 14056 19360 14062 19372
rect 14093 19363 14151 19369
rect 14093 19360 14105 19363
rect 14056 19332 14105 19360
rect 14056 19320 14062 19332
rect 14093 19329 14105 19332
rect 14139 19360 14151 19363
rect 14277 19363 14335 19369
rect 14277 19360 14289 19363
rect 14139 19332 14289 19360
rect 14139 19329 14151 19332
rect 14093 19323 14151 19329
rect 14277 19329 14289 19332
rect 14323 19329 14335 19363
rect 14277 19323 14335 19329
rect 14568 19332 14964 19360
rect 8128 19264 8708 19292
rect 4356 19224 4384 19252
rect 4982 19224 4988 19236
rect 4356 19196 4988 19224
rect 4816 19168 4844 19196
rect 4982 19184 4988 19196
rect 5040 19184 5046 19236
rect 6086 19184 6092 19236
rect 6144 19184 6150 19236
rect 7926 19184 7932 19236
rect 7984 19224 7990 19236
rect 8389 19227 8447 19233
rect 8389 19224 8401 19227
rect 7984 19196 8401 19224
rect 7984 19184 7990 19196
rect 8389 19193 8401 19196
rect 8435 19193 8447 19227
rect 8680 19224 8708 19264
rect 8754 19252 8760 19304
rect 8812 19252 8818 19304
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19261 8907 19295
rect 8849 19255 8907 19261
rect 9033 19295 9091 19301
rect 9033 19261 9045 19295
rect 9079 19292 9091 19295
rect 9674 19292 9680 19304
rect 9079 19264 9680 19292
rect 9079 19261 9091 19264
rect 9033 19255 9091 19261
rect 8864 19224 8892 19255
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 10226 19252 10232 19304
rect 10284 19292 10290 19304
rect 10870 19292 10876 19304
rect 10284 19264 10876 19292
rect 10284 19252 10290 19264
rect 10870 19252 10876 19264
rect 10928 19252 10934 19304
rect 10962 19252 10968 19304
rect 11020 19252 11026 19304
rect 11606 19252 11612 19304
rect 11664 19252 11670 19304
rect 12066 19252 12072 19304
rect 12124 19252 12130 19304
rect 12250 19252 12256 19304
rect 12308 19252 12314 19304
rect 12802 19252 12808 19304
rect 12860 19252 12866 19304
rect 13173 19295 13231 19301
rect 13173 19261 13185 19295
rect 13219 19261 13231 19295
rect 13173 19255 13231 19261
rect 8680 19196 8892 19224
rect 8389 19187 8447 19193
rect 11698 19184 11704 19236
rect 11756 19224 11762 19236
rect 12268 19224 12296 19252
rect 11756 19196 12296 19224
rect 12820 19224 12848 19252
rect 13188 19224 13216 19255
rect 13538 19252 13544 19304
rect 13596 19292 13602 19304
rect 13725 19295 13783 19301
rect 13725 19292 13737 19295
rect 13596 19264 13737 19292
rect 13596 19252 13602 19264
rect 13725 19261 13737 19264
rect 13771 19261 13783 19295
rect 13725 19255 13783 19261
rect 14182 19252 14188 19304
rect 14240 19292 14246 19304
rect 14568 19292 14596 19332
rect 14936 19304 14964 19332
rect 14240 19264 14596 19292
rect 14240 19252 14246 19264
rect 14642 19252 14648 19304
rect 14700 19252 14706 19304
rect 14918 19252 14924 19304
rect 14976 19252 14982 19304
rect 15028 19292 15056 19400
rect 18141 19397 18153 19431
rect 18187 19397 18199 19431
rect 18141 19391 18199 19397
rect 16850 19320 16856 19372
rect 16908 19320 16914 19372
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19360 17371 19363
rect 18156 19360 18184 19391
rect 17359 19332 17908 19360
rect 18156 19332 18368 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 15194 19292 15200 19304
rect 15028 19264 15200 19292
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 16758 19252 16764 19304
rect 16816 19252 16822 19304
rect 16868 19292 16896 19320
rect 17880 19304 17908 19332
rect 17221 19295 17279 19301
rect 17221 19292 17233 19295
rect 16868 19264 17233 19292
rect 17221 19261 17233 19264
rect 17267 19261 17279 19295
rect 17221 19255 17279 19261
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 12820 19196 13216 19224
rect 11756 19184 11762 19196
rect 13814 19184 13820 19236
rect 13872 19224 13878 19236
rect 14737 19227 14795 19233
rect 14737 19224 14749 19227
rect 13872 19196 14749 19224
rect 13872 19184 13878 19196
rect 14737 19193 14749 19196
rect 14783 19193 14795 19227
rect 16776 19224 16804 19252
rect 17420 19224 17448 19255
rect 17862 19252 17868 19304
rect 17920 19252 17926 19304
rect 17954 19252 17960 19304
rect 18012 19252 18018 19304
rect 18138 19252 18144 19304
rect 18196 19252 18202 19304
rect 18230 19252 18236 19304
rect 18288 19252 18294 19304
rect 18340 19292 18368 19332
rect 18417 19295 18475 19301
rect 18417 19292 18429 19295
rect 18340 19264 18429 19292
rect 18417 19261 18429 19264
rect 18463 19292 18475 19295
rect 18693 19295 18751 19301
rect 18693 19292 18705 19295
rect 18463 19264 18705 19292
rect 18463 19261 18475 19264
rect 18417 19255 18475 19261
rect 18693 19261 18705 19264
rect 18739 19261 18751 19295
rect 18693 19255 18751 19261
rect 18874 19252 18880 19304
rect 18932 19252 18938 19304
rect 19150 19252 19156 19304
rect 19208 19252 19214 19304
rect 21082 19301 21088 19304
rect 20809 19295 20867 19301
rect 20809 19261 20821 19295
rect 20855 19261 20867 19295
rect 21076 19292 21088 19301
rect 21043 19264 21088 19292
rect 20809 19255 20867 19261
rect 21076 19255 21088 19264
rect 16776 19196 17448 19224
rect 19420 19227 19478 19233
rect 14737 19187 14795 19193
rect 19420 19193 19432 19227
rect 19466 19224 19478 19227
rect 19518 19224 19524 19236
rect 19466 19196 19524 19224
rect 19466 19193 19478 19196
rect 19420 19187 19478 19193
rect 19518 19184 19524 19196
rect 19576 19184 19582 19236
rect 20824 19224 20852 19255
rect 21082 19252 21088 19255
rect 21140 19252 21146 19304
rect 22465 19295 22523 19301
rect 22465 19292 22477 19295
rect 22066 19264 22477 19292
rect 21174 19224 21180 19236
rect 20824 19196 21180 19224
rect 21174 19184 21180 19196
rect 21232 19184 21238 19236
rect 4798 19116 4804 19168
rect 4856 19116 4862 19168
rect 5629 19159 5687 19165
rect 5629 19125 5641 19159
rect 5675 19156 5687 19159
rect 5902 19156 5908 19168
rect 5675 19128 5908 19156
rect 5675 19125 5687 19128
rect 5629 19119 5687 19125
rect 5902 19116 5908 19128
rect 5960 19116 5966 19168
rect 8205 19159 8263 19165
rect 8205 19125 8217 19159
rect 8251 19156 8263 19159
rect 10318 19156 10324 19168
rect 8251 19128 10324 19156
rect 8251 19125 8263 19128
rect 8205 19119 8263 19125
rect 10318 19116 10324 19128
rect 10376 19116 10382 19168
rect 12805 19159 12863 19165
rect 12805 19125 12817 19159
rect 12851 19156 12863 19159
rect 14182 19156 14188 19168
rect 12851 19128 14188 19156
rect 12851 19125 12863 19128
rect 12805 19119 12863 19125
rect 14182 19116 14188 19128
rect 14240 19116 14246 19168
rect 14553 19159 14611 19165
rect 14553 19125 14565 19159
rect 14599 19156 14611 19159
rect 15010 19156 15016 19168
rect 14599 19128 15016 19156
rect 14599 19125 14611 19128
rect 14553 19119 14611 19125
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 17126 19116 17132 19168
rect 17184 19116 17190 19168
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 18325 19159 18383 19165
rect 18325 19156 18337 19159
rect 18012 19128 18337 19156
rect 18012 19116 18018 19128
rect 18325 19125 18337 19128
rect 18371 19125 18383 19159
rect 18325 19119 18383 19125
rect 20346 19116 20352 19168
rect 20404 19156 20410 19168
rect 20533 19159 20591 19165
rect 20533 19156 20545 19159
rect 20404 19128 20545 19156
rect 20404 19116 20410 19128
rect 20533 19125 20545 19128
rect 20579 19125 20591 19159
rect 20533 19119 20591 19125
rect 20622 19116 20628 19168
rect 20680 19156 20686 19168
rect 22066 19156 22094 19264
rect 22465 19261 22477 19264
rect 22511 19261 22523 19295
rect 22465 19255 22523 19261
rect 22646 19252 22652 19304
rect 22704 19252 22710 19304
rect 22830 19252 22836 19304
rect 22888 19252 22894 19304
rect 22554 19184 22560 19236
rect 22612 19184 22618 19236
rect 20680 19128 22094 19156
rect 20680 19116 20686 19128
rect 22278 19116 22284 19168
rect 22336 19116 22342 19168
rect 552 19066 23368 19088
rect 552 19014 4322 19066
rect 4374 19014 4386 19066
rect 4438 19014 4450 19066
rect 4502 19014 4514 19066
rect 4566 19014 4578 19066
rect 4630 19014 23368 19066
rect 552 18992 23368 19014
rect 7466 18912 7472 18964
rect 7524 18912 7530 18964
rect 7926 18912 7932 18964
rect 7984 18912 7990 18964
rect 8018 18912 8024 18964
rect 8076 18952 8082 18964
rect 12713 18955 12771 18961
rect 8076 18924 10088 18952
rect 8076 18912 8082 18924
rect 5261 18887 5319 18893
rect 5261 18853 5273 18887
rect 5307 18884 5319 18887
rect 5626 18884 5632 18896
rect 5307 18856 5632 18884
rect 5307 18853 5319 18856
rect 5261 18847 5319 18853
rect 5626 18844 5632 18856
rect 5684 18884 5690 18896
rect 6822 18884 6828 18896
rect 5684 18856 6828 18884
rect 5684 18844 5690 18856
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 7484 18884 7512 18912
rect 8754 18884 8760 18896
rect 7484 18856 8760 18884
rect 8754 18844 8760 18856
rect 8812 18884 8818 18896
rect 8812 18856 8892 18884
rect 8812 18844 8818 18856
rect 5166 18776 5172 18828
rect 5224 18776 5230 18828
rect 5442 18776 5448 18828
rect 5500 18776 5506 18828
rect 5810 18776 5816 18828
rect 5868 18816 5874 18828
rect 6641 18819 6699 18825
rect 6641 18816 6653 18819
rect 5868 18788 6653 18816
rect 5868 18776 5874 18788
rect 5445 18683 5503 18689
rect 5445 18649 5457 18683
rect 5491 18680 5503 18683
rect 6086 18680 6092 18692
rect 5491 18652 6092 18680
rect 5491 18649 5503 18652
rect 5445 18643 5503 18649
rect 6086 18640 6092 18652
rect 6144 18640 6150 18692
rect 6472 18680 6500 18788
rect 6641 18785 6653 18788
rect 6687 18785 6699 18819
rect 7561 18819 7619 18825
rect 7561 18816 7573 18819
rect 6641 18779 6699 18785
rect 6748 18788 7573 18816
rect 6546 18708 6552 18760
rect 6604 18748 6610 18760
rect 6748 18748 6776 18788
rect 7561 18785 7573 18788
rect 7607 18785 7619 18819
rect 7561 18779 7619 18785
rect 7745 18819 7803 18825
rect 7745 18785 7757 18819
rect 7791 18785 7803 18819
rect 7745 18779 7803 18785
rect 6604 18720 6776 18748
rect 6604 18708 6610 18720
rect 6822 18708 6828 18760
rect 6880 18748 6886 18760
rect 7760 18748 7788 18779
rect 8478 18776 8484 18828
rect 8536 18776 8542 18828
rect 8864 18757 8892 18856
rect 9582 18844 9588 18896
rect 9640 18844 9646 18896
rect 10060 18884 10088 18924
rect 12713 18921 12725 18955
rect 12759 18952 12771 18955
rect 12802 18952 12808 18964
rect 12759 18924 12808 18952
rect 12759 18921 12771 18924
rect 12713 18915 12771 18921
rect 12802 18912 12808 18924
rect 12860 18912 12866 18964
rect 13357 18955 13415 18961
rect 13357 18921 13369 18955
rect 13403 18952 13415 18955
rect 14642 18952 14648 18964
rect 13403 18924 14648 18952
rect 13403 18921 13415 18924
rect 13357 18915 13415 18921
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 17678 18912 17684 18964
rect 17736 18952 17742 18964
rect 18049 18955 18107 18961
rect 18049 18952 18061 18955
rect 17736 18924 18061 18952
rect 17736 18912 17742 18924
rect 18049 18921 18061 18924
rect 18095 18952 18107 18955
rect 18874 18952 18880 18964
rect 18095 18924 18880 18952
rect 18095 18921 18107 18924
rect 18049 18915 18107 18921
rect 18874 18912 18880 18924
rect 18932 18912 18938 18964
rect 19978 18912 19984 18964
rect 20036 18912 20042 18964
rect 20625 18955 20683 18961
rect 20625 18921 20637 18955
rect 20671 18952 20683 18955
rect 21818 18952 21824 18964
rect 20671 18924 21824 18952
rect 20671 18921 20683 18924
rect 20625 18915 20683 18921
rect 21818 18912 21824 18924
rect 21876 18912 21882 18964
rect 22554 18912 22560 18964
rect 22612 18952 22618 18964
rect 22741 18955 22799 18961
rect 22741 18952 22753 18955
rect 22612 18924 22753 18952
rect 22612 18912 22618 18924
rect 22741 18921 22753 18924
rect 22787 18921 22799 18955
rect 22741 18915 22799 18921
rect 10962 18884 10968 18896
rect 10060 18856 10968 18884
rect 8941 18819 8999 18825
rect 8941 18785 8953 18819
rect 8987 18816 8999 18819
rect 9030 18816 9036 18828
rect 8987 18788 9036 18816
rect 8987 18785 8999 18788
rect 8941 18779 8999 18785
rect 9030 18776 9036 18788
rect 9088 18776 9094 18828
rect 10060 18825 10088 18856
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 12820 18884 12848 18912
rect 16209 18887 16267 18893
rect 16209 18884 16221 18887
rect 12820 18856 13308 18884
rect 9401 18819 9459 18825
rect 9401 18816 9413 18819
rect 9324 18788 9413 18816
rect 6880 18720 7788 18748
rect 8573 18751 8631 18757
rect 6880 18708 6886 18720
rect 8573 18717 8585 18751
rect 8619 18717 8631 18751
rect 8573 18711 8631 18717
rect 8849 18751 8907 18757
rect 8849 18717 8861 18751
rect 8895 18717 8907 18751
rect 8849 18711 8907 18717
rect 6914 18680 6920 18692
rect 6472 18652 6920 18680
rect 6914 18640 6920 18652
rect 6972 18640 6978 18692
rect 8110 18640 8116 18692
rect 8168 18640 8174 18692
rect 8588 18680 8616 18711
rect 9324 18689 9352 18788
rect 9401 18785 9413 18788
rect 9447 18785 9459 18819
rect 9401 18779 9459 18785
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18785 10103 18819
rect 10045 18779 10103 18785
rect 10410 18776 10416 18828
rect 10468 18776 10474 18828
rect 11333 18819 11391 18825
rect 11333 18816 11345 18819
rect 10520 18788 11345 18816
rect 10318 18708 10324 18760
rect 10376 18708 10382 18760
rect 9309 18683 9367 18689
rect 9309 18680 9321 18683
rect 8588 18652 9321 18680
rect 9309 18649 9321 18652
rect 9355 18649 9367 18683
rect 9858 18680 9864 18692
rect 9309 18643 9367 18649
rect 9416 18652 9864 18680
rect 7190 18572 7196 18624
rect 7248 18612 7254 18624
rect 9416 18612 9444 18652
rect 9858 18640 9864 18652
rect 9916 18640 9922 18692
rect 9950 18640 9956 18692
rect 10008 18680 10014 18692
rect 10520 18680 10548 18788
rect 11333 18785 11345 18788
rect 11379 18785 11391 18819
rect 11333 18779 11391 18785
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11572 18788 11805 18816
rect 11572 18776 11578 18788
rect 11793 18785 11805 18788
rect 11839 18816 11851 18819
rect 12158 18816 12164 18828
rect 11839 18788 12164 18816
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 12158 18776 12164 18788
rect 12216 18816 12222 18828
rect 12345 18819 12403 18825
rect 12345 18816 12357 18819
rect 12216 18788 12357 18816
rect 12216 18776 12222 18788
rect 12345 18785 12357 18788
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 13078 18776 13084 18828
rect 13136 18776 13142 18828
rect 10870 18708 10876 18760
rect 10928 18748 10934 18760
rect 11057 18751 11115 18757
rect 11057 18748 11069 18751
rect 10928 18720 11069 18748
rect 10928 18708 10934 18720
rect 11057 18717 11069 18720
rect 11103 18717 11115 18751
rect 11974 18748 11980 18760
rect 11057 18711 11115 18717
rect 11716 18720 11980 18748
rect 10008 18652 10548 18680
rect 10781 18683 10839 18689
rect 10008 18640 10014 18652
rect 10781 18649 10793 18683
rect 10827 18680 10839 18683
rect 11716 18680 11744 18720
rect 11974 18708 11980 18720
rect 12032 18748 12038 18760
rect 12253 18751 12311 18757
rect 12253 18748 12265 18751
rect 12032 18720 12265 18748
rect 12032 18708 12038 18720
rect 12253 18717 12265 18720
rect 12299 18717 12311 18751
rect 12253 18711 12311 18717
rect 12986 18708 12992 18760
rect 13044 18748 13050 18760
rect 13173 18751 13231 18757
rect 13173 18748 13185 18751
rect 13044 18720 13185 18748
rect 13044 18708 13050 18720
rect 13173 18717 13185 18720
rect 13219 18717 13231 18751
rect 13280 18748 13308 18856
rect 13464 18856 16221 18884
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 13280 18720 13369 18748
rect 13173 18711 13231 18717
rect 13357 18717 13369 18720
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 10827 18652 11744 18680
rect 10827 18649 10839 18652
rect 10781 18643 10839 18649
rect 11790 18640 11796 18692
rect 11848 18680 11854 18692
rect 13464 18680 13492 18856
rect 13725 18819 13783 18825
rect 13725 18785 13737 18819
rect 13771 18816 13783 18819
rect 13814 18816 13820 18828
rect 13771 18788 13820 18816
rect 13771 18785 13783 18788
rect 13725 18779 13783 18785
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 14274 18776 14280 18828
rect 14332 18776 14338 18828
rect 14550 18776 14556 18828
rect 14608 18816 14614 18828
rect 14921 18819 14979 18825
rect 14921 18816 14933 18819
rect 14608 18788 14933 18816
rect 14608 18776 14614 18788
rect 14921 18785 14933 18788
rect 14967 18816 14979 18819
rect 15102 18816 15108 18828
rect 14967 18788 15108 18816
rect 14967 18785 14979 18788
rect 14921 18779 14979 18785
rect 15102 18776 15108 18788
rect 15160 18776 15166 18828
rect 15764 18825 15792 18856
rect 16209 18853 16221 18856
rect 16255 18884 16267 18887
rect 16758 18884 16764 18896
rect 16255 18856 16764 18884
rect 16255 18853 16267 18856
rect 16209 18847 16267 18853
rect 16758 18844 16764 18856
rect 16816 18844 16822 18896
rect 17126 18844 17132 18896
rect 17184 18884 17190 18896
rect 21628 18887 21686 18893
rect 17184 18856 17816 18884
rect 17184 18844 17190 18856
rect 15749 18819 15807 18825
rect 15749 18785 15761 18819
rect 15795 18785 15807 18819
rect 16117 18819 16175 18825
rect 16117 18816 16129 18819
rect 15749 18779 15807 18785
rect 15856 18788 16129 18816
rect 13998 18708 14004 18760
rect 14056 18708 14062 18760
rect 15856 18757 15884 18788
rect 16117 18785 16129 18788
rect 16163 18785 16175 18819
rect 16117 18779 16175 18785
rect 16390 18776 16396 18828
rect 16448 18776 16454 18828
rect 17788 18825 17816 18856
rect 21628 18853 21640 18887
rect 21674 18884 21686 18887
rect 22278 18884 22284 18896
rect 21674 18856 22284 18884
rect 21674 18853 21686 18856
rect 21628 18847 21686 18853
rect 22278 18844 22284 18856
rect 22336 18844 22342 18896
rect 17681 18819 17739 18825
rect 17681 18785 17693 18819
rect 17727 18785 17739 18819
rect 17681 18779 17739 18785
rect 17773 18819 17831 18825
rect 17773 18785 17785 18819
rect 17819 18816 17831 18819
rect 17957 18819 18015 18825
rect 17957 18816 17969 18819
rect 17819 18788 17969 18816
rect 17819 18785 17831 18788
rect 17773 18779 17831 18785
rect 17957 18785 17969 18788
rect 18003 18785 18015 18819
rect 17957 18779 18015 18785
rect 18141 18819 18199 18825
rect 18141 18785 18153 18819
rect 18187 18785 18199 18819
rect 18141 18779 18199 18785
rect 14185 18751 14243 18757
rect 14185 18717 14197 18751
rect 14231 18717 14243 18751
rect 14829 18751 14887 18757
rect 14829 18748 14841 18751
rect 14185 18711 14243 18717
rect 14292 18720 14841 18748
rect 11848 18652 13492 18680
rect 13541 18683 13599 18689
rect 11848 18640 11854 18652
rect 13541 18649 13553 18683
rect 13587 18680 13599 18683
rect 14200 18680 14228 18711
rect 13587 18652 14228 18680
rect 13587 18649 13599 18652
rect 13541 18643 13599 18649
rect 7248 18584 9444 18612
rect 7248 18572 7254 18584
rect 9766 18572 9772 18624
rect 9824 18572 9830 18624
rect 13906 18572 13912 18624
rect 13964 18572 13970 18624
rect 14182 18572 14188 18624
rect 14240 18612 14246 18624
rect 14292 18612 14320 18720
rect 14829 18717 14841 18720
rect 14875 18717 14887 18751
rect 14829 18711 14887 18717
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18748 15347 18751
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 15335 18720 15853 18748
rect 15335 18717 15347 18720
rect 15289 18711 15347 18717
rect 15841 18717 15853 18720
rect 15887 18717 15899 18751
rect 17696 18748 17724 18779
rect 18156 18748 18184 18779
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 20165 18819 20223 18825
rect 20165 18816 20177 18819
rect 19760 18788 20177 18816
rect 19760 18776 19766 18788
rect 20165 18785 20177 18788
rect 20211 18785 20223 18819
rect 20165 18779 20223 18785
rect 15841 18711 15899 18717
rect 16408 18720 18184 18748
rect 20180 18748 20208 18779
rect 20346 18776 20352 18828
rect 20404 18776 20410 18828
rect 20533 18819 20591 18825
rect 20533 18785 20545 18819
rect 20579 18816 20591 18819
rect 20622 18816 20628 18828
rect 20579 18788 20628 18816
rect 20579 18785 20591 18788
rect 20533 18779 20591 18785
rect 20548 18748 20576 18779
rect 20622 18776 20628 18788
rect 20680 18776 20686 18828
rect 21082 18776 21088 18828
rect 21140 18776 21146 18828
rect 22370 18776 22376 18828
rect 22428 18816 22434 18828
rect 22922 18816 22928 18828
rect 22428 18788 22928 18816
rect 22428 18776 22434 18788
rect 22922 18776 22928 18788
rect 22980 18816 22986 18828
rect 23017 18819 23075 18825
rect 23017 18816 23029 18819
rect 22980 18788 23029 18816
rect 22980 18776 22986 18788
rect 23017 18785 23029 18788
rect 23063 18785 23075 18819
rect 23017 18779 23075 18785
rect 20180 18720 20576 18748
rect 16408 18689 16436 18720
rect 16393 18683 16451 18689
rect 16393 18649 16405 18683
rect 16439 18649 16451 18683
rect 20548 18680 20576 18720
rect 21174 18708 21180 18760
rect 21232 18748 21238 18760
rect 21361 18751 21419 18757
rect 21361 18748 21373 18751
rect 21232 18720 21373 18748
rect 21232 18708 21238 18720
rect 21361 18717 21373 18720
rect 21407 18717 21419 18751
rect 21361 18711 21419 18717
rect 20901 18683 20959 18689
rect 20901 18680 20913 18683
rect 20548 18652 20913 18680
rect 16393 18643 16451 18649
rect 20901 18649 20913 18652
rect 20947 18649 20959 18683
rect 20901 18643 20959 18649
rect 14240 18584 14320 18612
rect 14553 18615 14611 18621
rect 14240 18572 14246 18584
rect 14553 18581 14565 18615
rect 14599 18612 14611 18615
rect 15286 18612 15292 18624
rect 14599 18584 15292 18612
rect 14599 18581 14611 18584
rect 14553 18575 14611 18581
rect 15286 18572 15292 18584
rect 15344 18572 15350 18624
rect 15470 18572 15476 18624
rect 15528 18612 15534 18624
rect 16482 18612 16488 18624
rect 15528 18584 16488 18612
rect 15528 18572 15534 18584
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 17497 18615 17555 18621
rect 17497 18581 17509 18615
rect 17543 18612 17555 18615
rect 17586 18612 17592 18624
rect 17543 18584 17592 18612
rect 17543 18581 17555 18584
rect 17497 18575 17555 18581
rect 17586 18572 17592 18584
rect 17644 18572 17650 18624
rect 21358 18572 21364 18624
rect 21416 18612 21422 18624
rect 22462 18612 22468 18624
rect 21416 18584 22468 18612
rect 21416 18572 21422 18584
rect 22462 18572 22468 18584
rect 22520 18572 22526 18624
rect 22925 18615 22983 18621
rect 22925 18581 22937 18615
rect 22971 18612 22983 18615
rect 23014 18612 23020 18624
rect 22971 18584 23020 18612
rect 22971 18581 22983 18584
rect 22925 18575 22983 18581
rect 23014 18572 23020 18584
rect 23072 18572 23078 18624
rect 552 18522 23368 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 23368 18522
rect 552 18448 23368 18470
rect 5353 18411 5411 18417
rect 5353 18377 5365 18411
rect 5399 18408 5411 18411
rect 6546 18408 6552 18420
rect 5399 18380 6552 18408
rect 5399 18377 5411 18380
rect 5353 18371 5411 18377
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 7101 18411 7159 18417
rect 7101 18377 7113 18411
rect 7147 18408 7159 18411
rect 14182 18408 14188 18420
rect 7147 18380 14188 18408
rect 7147 18377 7159 18380
rect 7101 18371 7159 18377
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 14274 18368 14280 18420
rect 14332 18408 14338 18420
rect 14921 18411 14979 18417
rect 14921 18408 14933 18411
rect 14332 18380 14933 18408
rect 14332 18368 14338 18380
rect 14921 18377 14933 18380
rect 14967 18377 14979 18411
rect 14921 18371 14979 18377
rect 15565 18411 15623 18417
rect 15565 18377 15577 18411
rect 15611 18408 15623 18411
rect 16390 18408 16396 18420
rect 15611 18380 16396 18408
rect 15611 18377 15623 18380
rect 15565 18371 15623 18377
rect 16390 18368 16396 18380
rect 16448 18368 16454 18420
rect 17773 18411 17831 18417
rect 17773 18377 17785 18411
rect 17819 18408 17831 18411
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 17819 18380 18061 18408
rect 17819 18377 17831 18380
rect 17773 18371 17831 18377
rect 18049 18377 18061 18380
rect 18095 18408 18107 18411
rect 18414 18408 18420 18420
rect 18095 18380 18420 18408
rect 18095 18377 18107 18380
rect 18049 18371 18107 18377
rect 18414 18368 18420 18380
rect 18472 18408 18478 18420
rect 21545 18411 21603 18417
rect 18472 18380 19012 18408
rect 18472 18368 18478 18380
rect 4617 18343 4675 18349
rect 4617 18309 4629 18343
rect 4663 18340 4675 18343
rect 5166 18340 5172 18352
rect 4663 18312 5172 18340
rect 4663 18309 4675 18312
rect 4617 18303 4675 18309
rect 5166 18300 5172 18312
rect 5224 18340 5230 18352
rect 8754 18340 8760 18352
rect 5224 18312 5580 18340
rect 5224 18300 5230 18312
rect 4154 18272 4160 18284
rect 4080 18244 4160 18272
rect 4080 18213 4108 18244
rect 4154 18232 4160 18244
rect 4212 18272 4218 18284
rect 4982 18272 4988 18284
rect 4212 18244 4988 18272
rect 4212 18232 4218 18244
rect 4982 18232 4988 18244
rect 5040 18272 5046 18284
rect 5552 18281 5580 18312
rect 8680 18312 8760 18340
rect 5537 18275 5595 18281
rect 5040 18244 5212 18272
rect 5040 18232 5046 18244
rect 4065 18207 4123 18213
rect 4065 18173 4077 18207
rect 4111 18173 4123 18207
rect 4065 18167 4123 18173
rect 4433 18207 4491 18213
rect 4433 18173 4445 18207
rect 4479 18204 4491 18207
rect 4614 18204 4620 18216
rect 4479 18176 4620 18204
rect 4479 18173 4491 18176
rect 4433 18167 4491 18173
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 4709 18207 4767 18213
rect 4709 18173 4721 18207
rect 4755 18204 4767 18207
rect 4755 18176 4789 18204
rect 4755 18173 4767 18176
rect 4709 18167 4767 18173
rect 4246 18096 4252 18148
rect 4304 18096 4310 18148
rect 4338 18096 4344 18148
rect 4396 18136 4402 18148
rect 4724 18136 4752 18167
rect 4890 18164 4896 18216
rect 4948 18164 4954 18216
rect 5184 18213 5212 18244
rect 5537 18241 5549 18275
rect 5583 18241 5595 18275
rect 5537 18235 5595 18241
rect 6181 18275 6239 18281
rect 6181 18241 6193 18275
rect 6227 18272 6239 18275
rect 6227 18244 6960 18272
rect 6227 18241 6239 18244
rect 6181 18235 6239 18241
rect 5169 18207 5227 18213
rect 5169 18173 5181 18207
rect 5215 18173 5227 18207
rect 5169 18167 5227 18173
rect 5626 18164 5632 18216
rect 5684 18164 5690 18216
rect 6086 18164 6092 18216
rect 6144 18164 6150 18216
rect 6932 18213 6960 18244
rect 6273 18207 6331 18213
rect 6273 18173 6285 18207
rect 6319 18173 6331 18207
rect 6273 18167 6331 18173
rect 6641 18207 6699 18213
rect 6641 18173 6653 18207
rect 6687 18173 6699 18207
rect 6641 18167 6699 18173
rect 6917 18207 6975 18213
rect 6917 18173 6929 18207
rect 6963 18173 6975 18207
rect 6917 18167 6975 18173
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 8680 18204 8708 18312
rect 8754 18300 8760 18312
rect 8812 18300 8818 18352
rect 9030 18300 9036 18352
rect 9088 18300 9094 18352
rect 14200 18340 14228 18368
rect 17589 18343 17647 18349
rect 14200 18312 15424 18340
rect 9048 18272 9076 18300
rect 8772 18244 9076 18272
rect 8772 18213 8800 18244
rect 10318 18232 10324 18284
rect 10376 18272 10382 18284
rect 10376 18244 11008 18272
rect 10376 18232 10382 18244
rect 8619 18176 8708 18204
rect 8757 18207 8815 18213
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 8757 18173 8769 18207
rect 8803 18173 8815 18207
rect 8757 18167 8815 18173
rect 8849 18207 8907 18213
rect 8849 18173 8861 18207
rect 8895 18173 8907 18207
rect 8849 18167 8907 18173
rect 9033 18207 9091 18213
rect 9033 18173 9045 18207
rect 9079 18204 9091 18207
rect 9306 18204 9312 18216
rect 9079 18176 9312 18204
rect 9079 18173 9091 18176
rect 9033 18167 9091 18173
rect 5074 18136 5080 18148
rect 4396 18108 5080 18136
rect 4396 18096 4402 18108
rect 5074 18096 5080 18108
rect 5132 18096 5138 18148
rect 6288 18136 6316 18167
rect 6012 18108 6316 18136
rect 6012 18080 6040 18108
rect 5994 18028 6000 18080
rect 6052 18028 6058 18080
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 6656 18068 6684 18167
rect 6733 18139 6791 18145
rect 6733 18105 6745 18139
rect 6779 18136 6791 18139
rect 7006 18136 7012 18148
rect 6779 18108 7012 18136
rect 6779 18105 6791 18108
rect 6733 18099 6791 18105
rect 7006 18096 7012 18108
rect 7064 18136 7070 18148
rect 7190 18136 7196 18148
rect 7064 18108 7196 18136
rect 7064 18096 7070 18108
rect 7190 18096 7196 18108
rect 7248 18096 7254 18148
rect 8478 18096 8484 18148
rect 8536 18136 8542 18148
rect 8864 18136 8892 18167
rect 9306 18164 9312 18176
rect 9364 18164 9370 18216
rect 10042 18164 10048 18216
rect 10100 18204 10106 18216
rect 10410 18204 10416 18216
rect 10100 18176 10416 18204
rect 10100 18164 10106 18176
rect 10410 18164 10416 18176
rect 10468 18204 10474 18216
rect 10980 18213 11008 18244
rect 11698 18232 11704 18284
rect 11756 18232 11762 18284
rect 11974 18232 11980 18284
rect 12032 18232 12038 18284
rect 13906 18232 13912 18284
rect 13964 18272 13970 18284
rect 14369 18275 14427 18281
rect 14369 18272 14381 18275
rect 13964 18244 14381 18272
rect 13964 18232 13970 18244
rect 14369 18241 14381 18244
rect 14415 18272 14427 18275
rect 14550 18272 14556 18284
rect 14415 18244 14556 18272
rect 14415 18241 14427 18244
rect 14369 18235 14427 18241
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 14642 18232 14648 18284
rect 14700 18232 14706 18284
rect 15102 18232 15108 18284
rect 15160 18272 15166 18284
rect 15197 18275 15255 18281
rect 15197 18272 15209 18275
rect 15160 18244 15209 18272
rect 15160 18232 15166 18244
rect 15197 18241 15209 18244
rect 15243 18241 15255 18275
rect 15197 18235 15255 18241
rect 10781 18207 10839 18213
rect 10781 18204 10793 18207
rect 10468 18176 10793 18204
rect 10468 18164 10474 18176
rect 10781 18173 10793 18176
rect 10827 18173 10839 18207
rect 10781 18167 10839 18173
rect 10965 18207 11023 18213
rect 10965 18173 10977 18207
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 11149 18207 11207 18213
rect 11149 18173 11161 18207
rect 11195 18204 11207 18207
rect 11241 18207 11299 18213
rect 11241 18204 11253 18207
rect 11195 18176 11253 18204
rect 11195 18173 11207 18176
rect 11149 18167 11207 18173
rect 11241 18173 11253 18176
rect 11287 18173 11299 18207
rect 11241 18167 11299 18173
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 12066 18204 12072 18216
rect 11931 18176 12072 18204
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 12066 18164 12072 18176
rect 12124 18164 12130 18216
rect 13998 18164 14004 18216
rect 14056 18204 14062 18216
rect 14277 18207 14335 18213
rect 14277 18204 14289 18207
rect 14056 18176 14289 18204
rect 14056 18164 14062 18176
rect 14277 18173 14289 18176
rect 14323 18173 14335 18207
rect 14277 18167 14335 18173
rect 14734 18164 14740 18216
rect 14792 18164 14798 18216
rect 14918 18164 14924 18216
rect 14976 18164 14982 18216
rect 15396 18213 15424 18312
rect 17589 18309 17601 18343
rect 17635 18340 17647 18343
rect 18138 18340 18144 18352
rect 17635 18312 18144 18340
rect 17635 18309 17647 18312
rect 17589 18303 17647 18309
rect 18138 18300 18144 18312
rect 18196 18340 18202 18352
rect 18984 18349 19012 18380
rect 21545 18377 21557 18411
rect 21591 18408 21603 18411
rect 21910 18408 21916 18420
rect 21591 18380 21916 18408
rect 21591 18377 21603 18380
rect 21545 18371 21603 18377
rect 21910 18368 21916 18380
rect 21968 18368 21974 18420
rect 22002 18368 22008 18420
rect 22060 18408 22066 18420
rect 22830 18408 22836 18420
rect 22060 18380 22836 18408
rect 22060 18368 22066 18380
rect 22830 18368 22836 18380
rect 22888 18368 22894 18420
rect 22922 18368 22928 18420
rect 22980 18408 22986 18420
rect 23017 18411 23075 18417
rect 23017 18408 23029 18411
rect 22980 18380 23029 18408
rect 22980 18368 22986 18380
rect 23017 18377 23029 18380
rect 23063 18377 23075 18411
rect 23017 18371 23075 18377
rect 18969 18343 19027 18349
rect 18196 18312 18460 18340
rect 18196 18300 18202 18312
rect 17420 18244 17724 18272
rect 17420 18213 17448 18244
rect 17696 18216 17724 18244
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18432 18281 18460 18312
rect 18969 18309 18981 18343
rect 19015 18309 19027 18343
rect 18969 18303 19027 18309
rect 18417 18275 18475 18281
rect 18012 18244 18368 18272
rect 18012 18232 18018 18244
rect 15381 18207 15439 18213
rect 15381 18173 15393 18207
rect 15427 18173 15439 18207
rect 15381 18167 15439 18173
rect 17405 18207 17463 18213
rect 17405 18173 17417 18207
rect 17451 18173 17463 18207
rect 17405 18167 17463 18173
rect 17586 18164 17592 18216
rect 17644 18164 17650 18216
rect 17678 18164 17684 18216
rect 17736 18164 17742 18216
rect 18230 18164 18236 18216
rect 18288 18164 18294 18216
rect 18340 18204 18368 18244
rect 18417 18241 18429 18275
rect 18463 18241 18475 18275
rect 18877 18275 18935 18281
rect 18877 18272 18889 18275
rect 18417 18235 18475 18241
rect 18524 18244 18889 18272
rect 18524 18204 18552 18244
rect 18877 18241 18889 18244
rect 18923 18241 18935 18275
rect 18877 18235 18935 18241
rect 21284 18244 21772 18272
rect 18340 18176 18552 18204
rect 18782 18164 18788 18216
rect 18840 18164 18846 18216
rect 18966 18164 18972 18216
rect 19024 18204 19030 18216
rect 19061 18207 19119 18213
rect 19061 18204 19073 18207
rect 19024 18176 19073 18204
rect 19024 18164 19030 18176
rect 19061 18173 19073 18176
rect 19107 18173 19119 18207
rect 19061 18167 19119 18173
rect 19245 18207 19303 18213
rect 19245 18173 19257 18207
rect 19291 18204 19303 18207
rect 19337 18207 19395 18213
rect 19337 18204 19349 18207
rect 19291 18176 19349 18204
rect 19291 18173 19303 18176
rect 19245 18167 19303 18173
rect 19337 18173 19349 18176
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 19702 18164 19708 18216
rect 19760 18164 19766 18216
rect 21284 18213 21312 18244
rect 21744 18216 21772 18244
rect 21269 18207 21327 18213
rect 21269 18173 21281 18207
rect 21315 18173 21327 18207
rect 21269 18167 21327 18173
rect 21358 18164 21364 18216
rect 21416 18204 21422 18216
rect 21637 18207 21695 18213
rect 21637 18204 21649 18207
rect 21416 18176 21649 18204
rect 21416 18164 21422 18176
rect 21637 18173 21649 18176
rect 21683 18173 21695 18207
rect 21637 18167 21695 18173
rect 21726 18164 21732 18216
rect 21784 18164 21790 18216
rect 22738 18204 22744 18216
rect 21836 18176 22744 18204
rect 9490 18136 9496 18148
rect 8536 18108 9496 18136
rect 8536 18096 8542 18108
rect 9490 18096 9496 18108
rect 9548 18096 9554 18148
rect 11425 18139 11483 18145
rect 11425 18105 11437 18139
rect 11471 18136 11483 18139
rect 12894 18136 12900 18148
rect 11471 18108 12900 18136
rect 11471 18105 11483 18108
rect 11425 18099 11483 18105
rect 12894 18096 12900 18108
rect 12952 18096 12958 18148
rect 17957 18139 18015 18145
rect 17957 18105 17969 18139
rect 18003 18136 18015 18139
rect 19521 18139 19579 18145
rect 19521 18136 19533 18139
rect 18003 18108 19533 18136
rect 18003 18105 18015 18108
rect 17957 18099 18015 18105
rect 19521 18105 19533 18108
rect 19567 18105 19579 18139
rect 19521 18099 19579 18105
rect 19613 18139 19671 18145
rect 19613 18105 19625 18139
rect 19659 18105 19671 18139
rect 19613 18099 19671 18105
rect 21545 18139 21603 18145
rect 21545 18105 21557 18139
rect 21591 18136 21603 18139
rect 21836 18136 21864 18176
rect 22738 18164 22744 18176
rect 22796 18164 22802 18216
rect 21910 18145 21916 18148
rect 21591 18108 21864 18136
rect 21591 18105 21603 18108
rect 21545 18099 21603 18105
rect 21904 18099 21916 18145
rect 21968 18136 21974 18148
rect 21968 18108 22004 18136
rect 6328 18040 6684 18068
rect 6328 18028 6334 18040
rect 8754 18028 8760 18080
rect 8812 18028 8818 18080
rect 8846 18028 8852 18080
rect 8904 18028 8910 18080
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 19628 18068 19656 18099
rect 21910 18096 21916 18099
rect 21968 18096 21974 18108
rect 18656 18040 19656 18068
rect 18656 18028 18662 18040
rect 19886 18028 19892 18080
rect 19944 18028 19950 18080
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 22922 18068 22928 18080
rect 21407 18040 22928 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 22922 18028 22928 18040
rect 22980 18028 22986 18080
rect 552 17978 23368 18000
rect 552 17926 4322 17978
rect 4374 17926 4386 17978
rect 4438 17926 4450 17978
rect 4502 17926 4514 17978
rect 4566 17926 4578 17978
rect 4630 17926 23368 17978
rect 552 17904 23368 17926
rect 4065 17867 4123 17873
rect 4065 17833 4077 17867
rect 4111 17864 4123 17867
rect 4154 17864 4160 17876
rect 4111 17836 4160 17864
rect 4111 17833 4123 17836
rect 4065 17827 4123 17833
rect 4154 17824 4160 17836
rect 4212 17824 4218 17876
rect 8754 17824 8760 17876
rect 8812 17864 8818 17876
rect 9125 17867 9183 17873
rect 9125 17864 9137 17867
rect 8812 17836 9137 17864
rect 8812 17824 8818 17836
rect 9125 17833 9137 17836
rect 9171 17864 9183 17867
rect 9398 17864 9404 17876
rect 9171 17836 9404 17864
rect 9171 17833 9183 17836
rect 9125 17827 9183 17833
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 10042 17824 10048 17876
rect 10100 17824 10106 17876
rect 18233 17867 18291 17873
rect 18233 17833 18245 17867
rect 18279 17864 18291 17867
rect 18506 17864 18512 17876
rect 18279 17836 18512 17864
rect 18279 17833 18291 17836
rect 18233 17827 18291 17833
rect 18506 17824 18512 17836
rect 18564 17824 18570 17876
rect 18598 17824 18604 17876
rect 18656 17824 18662 17876
rect 22738 17824 22744 17876
rect 22796 17824 22802 17876
rect 3789 17799 3847 17805
rect 3789 17765 3801 17799
rect 3835 17796 3847 17799
rect 4798 17796 4804 17808
rect 3835 17768 4804 17796
rect 3835 17765 3847 17768
rect 3789 17759 3847 17765
rect 4632 17740 4660 17768
rect 4798 17756 4804 17768
rect 4856 17756 4862 17808
rect 5626 17796 5632 17808
rect 5184 17768 5632 17796
rect 4338 17688 4344 17740
rect 4396 17688 4402 17740
rect 4614 17688 4620 17740
rect 4672 17688 4678 17740
rect 5184 17737 5212 17768
rect 5626 17756 5632 17768
rect 5684 17796 5690 17808
rect 9766 17796 9772 17808
rect 5684 17768 6132 17796
rect 5684 17756 5690 17768
rect 5169 17731 5227 17737
rect 5169 17697 5181 17731
rect 5215 17697 5227 17731
rect 5902 17728 5908 17740
rect 5169 17691 5227 17697
rect 5276 17700 5908 17728
rect 4430 17620 4436 17672
rect 4488 17660 4494 17672
rect 4890 17660 4896 17672
rect 4488 17632 4896 17660
rect 4488 17620 4494 17632
rect 4890 17620 4896 17632
rect 4948 17620 4954 17672
rect 4985 17663 5043 17669
rect 4985 17629 4997 17663
rect 5031 17660 5043 17663
rect 5276 17660 5304 17700
rect 5902 17688 5908 17700
rect 5960 17688 5966 17740
rect 6104 17737 6132 17768
rect 9048 17768 9772 17796
rect 6089 17731 6147 17737
rect 6089 17697 6101 17731
rect 6135 17697 6147 17731
rect 6089 17691 6147 17697
rect 6917 17731 6975 17737
rect 6917 17697 6929 17731
rect 6963 17728 6975 17731
rect 7374 17728 7380 17740
rect 6963 17700 7380 17728
rect 6963 17697 6975 17700
rect 6917 17691 6975 17697
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 7466 17688 7472 17740
rect 7524 17728 7530 17740
rect 9048 17737 9076 17768
rect 9766 17756 9772 17768
rect 9824 17756 9830 17808
rect 13906 17756 13912 17808
rect 13964 17796 13970 17808
rect 19736 17799 19794 17805
rect 13964 17768 16620 17796
rect 13964 17756 13970 17768
rect 7561 17731 7619 17737
rect 7561 17728 7573 17731
rect 7524 17700 7573 17728
rect 7524 17688 7530 17700
rect 7561 17697 7573 17700
rect 7607 17697 7619 17731
rect 7561 17691 7619 17697
rect 9033 17731 9091 17737
rect 9033 17697 9045 17731
rect 9079 17697 9091 17731
rect 9033 17691 9091 17697
rect 9309 17731 9367 17737
rect 9309 17697 9321 17731
rect 9355 17728 9367 17731
rect 9490 17728 9496 17740
rect 9355 17700 9496 17728
rect 9355 17697 9367 17700
rect 9309 17691 9367 17697
rect 9490 17688 9496 17700
rect 9548 17688 9554 17740
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17697 9735 17731
rect 9677 17691 9735 17697
rect 5031 17632 5304 17660
rect 5537 17663 5595 17669
rect 5031 17629 5043 17632
rect 4985 17623 5043 17629
rect 5537 17629 5549 17663
rect 5583 17660 5595 17663
rect 5626 17660 5632 17672
rect 5583 17632 5632 17660
rect 5583 17629 5595 17632
rect 5537 17623 5595 17629
rect 5626 17620 5632 17632
rect 5684 17620 5690 17672
rect 5445 17595 5503 17601
rect 5445 17561 5457 17595
rect 5491 17592 5503 17595
rect 6086 17592 6092 17604
rect 5491 17564 6092 17592
rect 5491 17561 5503 17564
rect 5445 17555 5503 17561
rect 6086 17552 6092 17564
rect 6144 17552 6150 17604
rect 9214 17552 9220 17604
rect 9272 17592 9278 17604
rect 9692 17592 9720 17691
rect 14918 17688 14924 17740
rect 14976 17728 14982 17740
rect 16301 17731 16359 17737
rect 16301 17728 16313 17731
rect 14976 17700 16313 17728
rect 14976 17688 14982 17700
rect 16301 17697 16313 17700
rect 16347 17697 16359 17731
rect 16301 17691 16359 17697
rect 9769 17663 9827 17669
rect 9769 17629 9781 17663
rect 9815 17660 9827 17663
rect 9858 17660 9864 17672
rect 9815 17632 9864 17660
rect 9815 17629 9827 17632
rect 9769 17623 9827 17629
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 16316 17660 16344 17691
rect 16482 17688 16488 17740
rect 16540 17688 16546 17740
rect 16592 17737 16620 17768
rect 19736 17765 19748 17799
rect 19782 17796 19794 17799
rect 19886 17796 19892 17808
rect 19782 17768 19892 17796
rect 19782 17765 19794 17768
rect 19736 17759 19794 17765
rect 19886 17756 19892 17768
rect 19944 17756 19950 17808
rect 21085 17799 21143 17805
rect 21085 17765 21097 17799
rect 21131 17796 21143 17799
rect 21514 17799 21572 17805
rect 21514 17796 21526 17799
rect 21131 17768 21526 17796
rect 21131 17765 21143 17768
rect 21085 17759 21143 17765
rect 21514 17765 21526 17768
rect 21560 17765 21572 17799
rect 21514 17759 21572 17765
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 16666 17728 16672 17740
rect 16623 17700 16672 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 16666 17688 16672 17700
rect 16724 17688 16730 17740
rect 17218 17688 17224 17740
rect 17276 17688 17282 17740
rect 17405 17731 17463 17737
rect 17405 17697 17417 17731
rect 17451 17697 17463 17731
rect 17405 17691 17463 17697
rect 16850 17660 16856 17672
rect 16316 17632 16856 17660
rect 16850 17620 16856 17632
rect 16908 17620 16914 17672
rect 17420 17660 17448 17691
rect 17586 17688 17592 17740
rect 17644 17688 17650 17740
rect 17865 17731 17923 17737
rect 17865 17697 17877 17731
rect 17911 17728 17923 17731
rect 17954 17728 17960 17740
rect 17911 17700 17960 17728
rect 17911 17697 17923 17700
rect 17865 17691 17923 17697
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 18138 17688 18144 17740
rect 18196 17688 18202 17740
rect 18230 17688 18236 17740
rect 18288 17728 18294 17740
rect 18325 17731 18383 17737
rect 18325 17728 18337 17731
rect 18288 17700 18337 17728
rect 18288 17688 18294 17700
rect 18325 17697 18337 17700
rect 18371 17697 18383 17731
rect 18325 17691 18383 17697
rect 18509 17731 18567 17737
rect 18509 17697 18521 17731
rect 18555 17697 18567 17731
rect 18509 17691 18567 17697
rect 17144 17632 17448 17660
rect 18156 17660 18184 17688
rect 18524 17660 18552 17691
rect 18690 17688 18696 17740
rect 18748 17728 18754 17740
rect 19150 17728 19156 17740
rect 18748 17700 19156 17728
rect 18748 17688 18754 17700
rect 19150 17688 19156 17700
rect 19208 17728 19214 17740
rect 19981 17731 20039 17737
rect 19981 17728 19993 17731
rect 19208 17700 19993 17728
rect 19208 17688 19214 17700
rect 19981 17697 19993 17700
rect 20027 17728 20039 17731
rect 20027 17700 20760 17728
rect 20027 17697 20039 17700
rect 19981 17691 20039 17697
rect 18156 17632 18552 17660
rect 20625 17663 20683 17669
rect 17144 17604 17172 17632
rect 20625 17629 20637 17663
rect 20671 17629 20683 17663
rect 20732 17660 20760 17700
rect 20898 17688 20904 17740
rect 20956 17688 20962 17740
rect 22002 17688 22008 17740
rect 22060 17728 22066 17740
rect 22060 17700 22784 17728
rect 22060 17688 22066 17700
rect 21174 17660 21180 17672
rect 20732 17632 21180 17660
rect 20625 17623 20683 17629
rect 9272 17564 9720 17592
rect 9272 17552 9278 17564
rect 17126 17552 17132 17604
rect 17184 17552 17190 17604
rect 20640 17592 20668 17623
rect 21174 17620 21180 17632
rect 21232 17660 21238 17672
rect 22756 17669 22784 17700
rect 22830 17688 22836 17740
rect 22888 17728 22894 17740
rect 22925 17731 22983 17737
rect 22925 17728 22937 17731
rect 22888 17700 22937 17728
rect 22888 17688 22894 17700
rect 22925 17697 22937 17700
rect 22971 17697 22983 17731
rect 22925 17691 22983 17697
rect 23014 17688 23020 17740
rect 23072 17688 23078 17740
rect 21269 17663 21327 17669
rect 21269 17660 21281 17663
rect 21232 17632 21281 17660
rect 21232 17620 21238 17632
rect 21269 17629 21281 17632
rect 21315 17629 21327 17663
rect 21269 17623 21327 17629
rect 22741 17663 22799 17669
rect 22741 17629 22753 17663
rect 22787 17629 22799 17663
rect 22741 17623 22799 17629
rect 20640 17564 21312 17592
rect 4706 17484 4712 17536
rect 4764 17484 4770 17536
rect 7561 17527 7619 17533
rect 7561 17493 7573 17527
rect 7607 17524 7619 17527
rect 8846 17524 8852 17536
rect 7607 17496 8852 17524
rect 7607 17493 7619 17496
rect 7561 17487 7619 17493
rect 8846 17484 8852 17496
rect 8904 17484 8910 17536
rect 9309 17527 9367 17533
rect 9309 17493 9321 17527
rect 9355 17524 9367 17527
rect 9858 17524 9864 17536
rect 9355 17496 9864 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 9858 17484 9864 17496
rect 9916 17484 9922 17536
rect 16117 17527 16175 17533
rect 16117 17493 16129 17527
rect 16163 17524 16175 17527
rect 16298 17524 16304 17536
rect 16163 17496 16304 17524
rect 16163 17493 16175 17496
rect 16117 17487 16175 17493
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 16669 17527 16727 17533
rect 16669 17493 16681 17527
rect 16715 17524 16727 17527
rect 16758 17524 16764 17536
rect 16715 17496 16764 17524
rect 16715 17493 16727 17496
rect 16669 17487 16727 17493
rect 16758 17484 16764 17496
rect 16816 17484 16822 17536
rect 18322 17484 18328 17536
rect 18380 17484 18386 17536
rect 18782 17484 18788 17536
rect 18840 17524 18846 17536
rect 20714 17524 20720 17536
rect 18840 17496 20720 17524
rect 18840 17484 18846 17496
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 21284 17524 21312 17564
rect 21542 17524 21548 17536
rect 21284 17496 21548 17524
rect 21542 17484 21548 17496
rect 21600 17524 21606 17536
rect 22649 17527 22707 17533
rect 22649 17524 22661 17527
rect 21600 17496 22661 17524
rect 21600 17484 21606 17496
rect 22649 17493 22661 17496
rect 22695 17493 22707 17527
rect 22649 17487 22707 17493
rect 552 17434 23368 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 23368 17434
rect 552 17360 23368 17382
rect 4246 17280 4252 17332
rect 4304 17320 4310 17332
rect 4525 17323 4583 17329
rect 4525 17320 4537 17323
rect 4304 17292 4537 17320
rect 4304 17280 4310 17292
rect 4525 17289 4537 17292
rect 4571 17289 4583 17323
rect 4525 17283 4583 17289
rect 4157 17119 4215 17125
rect 4157 17085 4169 17119
rect 4203 17116 4215 17119
rect 4430 17116 4436 17128
rect 4203 17088 4436 17116
rect 4203 17085 4215 17088
rect 4157 17079 4215 17085
rect 4430 17076 4436 17088
rect 4488 17076 4494 17128
rect 4540 17116 4568 17283
rect 4706 17280 4712 17332
rect 4764 17320 4770 17332
rect 5445 17323 5503 17329
rect 5445 17320 5457 17323
rect 4764 17292 5457 17320
rect 4764 17280 4770 17292
rect 5445 17289 5457 17292
rect 5491 17289 5503 17323
rect 5445 17283 5503 17289
rect 5626 17280 5632 17332
rect 5684 17280 5690 17332
rect 9490 17280 9496 17332
rect 9548 17280 9554 17332
rect 13906 17280 13912 17332
rect 13964 17280 13970 17332
rect 15933 17323 15991 17329
rect 15933 17289 15945 17323
rect 15979 17289 15991 17323
rect 15933 17283 15991 17289
rect 4985 17255 5043 17261
rect 4985 17221 4997 17255
rect 5031 17252 5043 17255
rect 7466 17252 7472 17264
rect 5031 17224 7472 17252
rect 5031 17221 5043 17224
rect 4985 17215 5043 17221
rect 5169 17187 5227 17193
rect 5169 17153 5181 17187
rect 5215 17184 5227 17187
rect 5534 17184 5540 17196
rect 5215 17156 5540 17184
rect 5215 17153 5227 17156
rect 5169 17147 5227 17153
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 5994 17144 6000 17196
rect 6052 17144 6058 17196
rect 6270 17144 6276 17196
rect 6328 17144 6334 17196
rect 7300 17193 7328 17224
rect 7466 17212 7472 17224
rect 7524 17212 7530 17264
rect 12529 17255 12587 17261
rect 12529 17221 12541 17255
rect 12575 17221 12587 17255
rect 12529 17215 12587 17221
rect 13357 17255 13415 17261
rect 13357 17221 13369 17255
rect 13403 17252 13415 17255
rect 15654 17252 15660 17264
rect 13403 17224 15660 17252
rect 13403 17221 13415 17224
rect 13357 17215 13415 17221
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17184 8263 17187
rect 9677 17187 9735 17193
rect 9677 17184 9689 17187
rect 8251 17156 9689 17184
rect 8251 17153 8263 17156
rect 8205 17147 8263 17153
rect 4617 17119 4675 17125
rect 4617 17116 4629 17119
rect 4540 17088 4629 17116
rect 4617 17085 4629 17088
rect 4663 17085 4675 17119
rect 4617 17079 4675 17085
rect 4982 17076 4988 17128
rect 5040 17076 5046 17128
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17116 5963 17119
rect 6086 17116 6092 17128
rect 5951 17088 6092 17116
rect 5951 17085 5963 17088
rect 5905 17079 5963 17085
rect 6086 17076 6092 17088
rect 6144 17076 6150 17128
rect 7374 17076 7380 17128
rect 7432 17076 7438 17128
rect 8846 17076 8852 17128
rect 8904 17076 8910 17128
rect 9140 17125 9168 17156
rect 9677 17153 9689 17156
rect 9723 17153 9735 17187
rect 9677 17147 9735 17153
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17184 10195 17187
rect 10597 17187 10655 17193
rect 10183 17156 10364 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 9125 17119 9183 17125
rect 9125 17085 9137 17119
rect 9171 17116 9183 17119
rect 9214 17116 9220 17128
rect 9171 17088 9220 17116
rect 9171 17085 9183 17088
rect 9125 17079 9183 17085
rect 9214 17076 9220 17088
rect 9272 17076 9278 17128
rect 9309 17119 9367 17125
rect 9309 17085 9321 17119
rect 9355 17116 9367 17119
rect 9769 17119 9827 17125
rect 9769 17116 9781 17119
rect 9355 17088 9781 17116
rect 9355 17085 9367 17088
rect 9309 17079 9367 17085
rect 9769 17085 9781 17088
rect 9815 17116 9827 17119
rect 9950 17116 9956 17128
rect 9815 17088 9956 17116
rect 9815 17085 9827 17088
rect 9769 17079 9827 17085
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 4338 17008 4344 17060
rect 4396 17048 4402 17060
rect 5074 17048 5080 17060
rect 4396 17020 5080 17048
rect 4396 17008 4402 17020
rect 5074 17008 5080 17020
rect 5132 17048 5138 17060
rect 5261 17051 5319 17057
rect 5261 17048 5273 17051
rect 5132 17020 5273 17048
rect 5132 17008 5138 17020
rect 5261 17017 5273 17020
rect 5307 17017 5319 17051
rect 5261 17011 5319 17017
rect 9030 17008 9036 17060
rect 9088 17048 9094 17060
rect 10152 17048 10180 17147
rect 10226 17076 10232 17128
rect 10284 17076 10290 17128
rect 10336 17116 10364 17156
rect 10597 17153 10609 17187
rect 10643 17184 10655 17187
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 10643 17156 11805 17184
rect 10643 17153 10655 17156
rect 10597 17147 10655 17153
rect 11793 17153 11805 17156
rect 11839 17184 11851 17187
rect 12069 17187 12127 17193
rect 12069 17184 12081 17187
rect 11839 17156 12081 17184
rect 11839 17153 11851 17156
rect 11793 17147 11851 17153
rect 12069 17153 12081 17156
rect 12115 17153 12127 17187
rect 12069 17147 12127 17153
rect 10689 17119 10747 17125
rect 10689 17118 10701 17119
rect 10612 17116 10701 17118
rect 10336 17090 10701 17116
rect 10336 17088 10640 17090
rect 10689 17085 10701 17090
rect 10735 17085 10747 17119
rect 10689 17079 10747 17085
rect 10870 17076 10876 17128
rect 10928 17076 10934 17128
rect 11698 17076 11704 17128
rect 11756 17116 11762 17128
rect 12161 17119 12219 17125
rect 12161 17116 12173 17119
rect 11756 17088 12173 17116
rect 11756 17076 11762 17088
rect 12161 17085 12173 17088
rect 12207 17085 12219 17119
rect 12544 17116 12572 17215
rect 15654 17212 15660 17224
rect 15712 17212 15718 17264
rect 15948 17252 15976 17283
rect 16482 17280 16488 17332
rect 16540 17320 16546 17332
rect 16540 17292 17080 17320
rect 16540 17280 16546 17292
rect 16853 17255 16911 17261
rect 16853 17252 16865 17255
rect 15948 17224 16865 17252
rect 12894 17144 12900 17196
rect 12952 17144 12958 17196
rect 14918 17184 14924 17196
rect 13832 17156 14924 17184
rect 12989 17119 13047 17125
rect 12989 17116 13001 17119
rect 12544 17088 13001 17116
rect 12161 17079 12219 17085
rect 12989 17085 13001 17088
rect 13035 17116 13047 17119
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 13035 17088 13737 17116
rect 13035 17085 13047 17088
rect 12989 17079 13047 17085
rect 13725 17085 13737 17088
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 9088 17020 10180 17048
rect 10781 17051 10839 17057
rect 9088 17008 9094 17020
rect 10781 17017 10793 17051
rect 10827 17048 10839 17051
rect 11149 17051 11207 17057
rect 11149 17048 11161 17051
rect 10827 17020 11161 17048
rect 10827 17017 10839 17020
rect 10781 17011 10839 17017
rect 11149 17017 11161 17020
rect 11195 17017 11207 17051
rect 11149 17011 11207 17017
rect 12894 17008 12900 17060
rect 12952 17048 12958 17060
rect 13541 17051 13599 17057
rect 13541 17048 13553 17051
rect 12952 17020 13553 17048
rect 12952 17008 12958 17020
rect 13541 17017 13553 17020
rect 13587 17017 13599 17051
rect 13541 17011 13599 17017
rect 4430 16940 4436 16992
rect 4488 16980 4494 16992
rect 5166 16980 5172 16992
rect 4488 16952 5172 16980
rect 4488 16940 4494 16952
rect 5166 16940 5172 16952
rect 5224 16980 5230 16992
rect 5461 16983 5519 16989
rect 5461 16980 5473 16983
rect 5224 16952 5473 16980
rect 5224 16940 5230 16952
rect 5461 16949 5473 16952
rect 5507 16949 5519 16983
rect 5461 16943 5519 16949
rect 8662 16940 8668 16992
rect 8720 16940 8726 16992
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 10870 16980 10876 16992
rect 10284 16952 10876 16980
rect 10284 16940 10290 16952
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 11701 16983 11759 16989
rect 11701 16949 11713 16983
rect 11747 16980 11759 16983
rect 13832 16980 13860 17156
rect 14918 17144 14924 17156
rect 14976 17144 14982 17196
rect 15749 17187 15807 17193
rect 15749 17153 15761 17187
rect 15795 17184 15807 17187
rect 15795 17156 16344 17184
rect 15795 17153 15807 17156
rect 15749 17147 15807 17153
rect 16316 17128 16344 17156
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17116 15071 17119
rect 15470 17116 15476 17128
rect 15059 17088 15476 17116
rect 15059 17085 15071 17088
rect 15013 17079 15071 17085
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 15654 17076 15660 17128
rect 15712 17116 15718 17128
rect 16025 17119 16083 17125
rect 16025 17116 16037 17119
rect 15712 17088 16037 17116
rect 15712 17076 15718 17088
rect 16025 17085 16037 17088
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 16298 17076 16304 17128
rect 16356 17076 16362 17128
rect 16592 17125 16620 17224
rect 16853 17221 16865 17224
rect 16899 17221 16911 17255
rect 16853 17215 16911 17221
rect 16577 17119 16635 17125
rect 16577 17085 16589 17119
rect 16623 17085 16635 17119
rect 16577 17079 16635 17085
rect 16758 17076 16764 17128
rect 16816 17076 16822 17128
rect 16850 17076 16856 17128
rect 16908 17076 16914 17128
rect 17052 17125 17080 17292
rect 17126 17280 17132 17332
rect 17184 17280 17190 17332
rect 17497 17323 17555 17329
rect 17497 17289 17509 17323
rect 17543 17320 17555 17323
rect 18230 17320 18236 17332
rect 17543 17292 18236 17320
rect 17543 17289 17555 17292
rect 17497 17283 17555 17289
rect 18230 17280 18236 17292
rect 18288 17280 18294 17332
rect 18322 17280 18328 17332
rect 18380 17280 18386 17332
rect 20898 17280 20904 17332
rect 20956 17320 20962 17332
rect 21082 17320 21088 17332
rect 20956 17292 21088 17320
rect 20956 17280 20962 17292
rect 21082 17280 21088 17292
rect 21140 17320 21146 17332
rect 22002 17320 22008 17332
rect 21140 17292 22008 17320
rect 21140 17280 21146 17292
rect 22002 17280 22008 17292
rect 22060 17320 22066 17332
rect 22373 17323 22431 17329
rect 22373 17320 22385 17323
rect 22060 17292 22385 17320
rect 22060 17280 22066 17292
rect 22373 17289 22385 17292
rect 22419 17289 22431 17323
rect 22373 17283 22431 17289
rect 17586 17184 17592 17196
rect 17144 17156 17592 17184
rect 17144 17125 17172 17156
rect 17586 17144 17592 17156
rect 17644 17144 17650 17196
rect 18187 17187 18245 17193
rect 18187 17153 18199 17187
rect 18233 17184 18245 17187
rect 18414 17184 18420 17196
rect 18233 17156 18420 17184
rect 18233 17153 18245 17156
rect 18187 17147 18245 17153
rect 18414 17144 18420 17156
rect 18472 17144 18478 17196
rect 17037 17119 17095 17125
rect 17037 17085 17049 17119
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 16117 17051 16175 17057
rect 16117 17017 16129 17051
rect 16163 17048 16175 17051
rect 17144 17048 17172 17079
rect 17218 17076 17224 17128
rect 17276 17076 17282 17128
rect 18046 17076 18052 17128
rect 18104 17076 18110 17128
rect 18506 17076 18512 17128
rect 18564 17076 18570 17128
rect 18690 17076 18696 17128
rect 18748 17076 18754 17128
rect 16163 17020 17172 17048
rect 16163 17017 16175 17020
rect 16117 17011 16175 17017
rect 11747 16952 13860 16980
rect 11747 16949 11759 16952
rect 11701 16943 11759 16949
rect 15378 16940 15384 16992
rect 15436 16940 15442 16992
rect 15473 16983 15531 16989
rect 15473 16949 15485 16983
rect 15519 16980 15531 16983
rect 15562 16980 15568 16992
rect 15519 16952 15568 16980
rect 15519 16949 15531 16952
rect 15473 16943 15531 16949
rect 15562 16940 15568 16952
rect 15620 16940 15626 16992
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 17236 16980 17264 17076
rect 18417 17051 18475 17057
rect 18417 17017 18429 17051
rect 18463 17048 18475 17051
rect 18938 17051 18996 17057
rect 18938 17048 18950 17051
rect 18463 17020 18950 17048
rect 18463 17017 18475 17020
rect 18417 17011 18475 17017
rect 18938 17017 18950 17020
rect 18984 17017 18996 17051
rect 18938 17011 18996 17017
rect 22649 17051 22707 17057
rect 22649 17017 22661 17051
rect 22695 17048 22707 17051
rect 22738 17048 22744 17060
rect 22695 17020 22744 17048
rect 22695 17017 22707 17020
rect 22649 17011 22707 17017
rect 22738 17008 22744 17020
rect 22796 17008 22802 17060
rect 16080 16952 17264 16980
rect 16080 16940 16086 16952
rect 19242 16940 19248 16992
rect 19300 16980 19306 16992
rect 20073 16983 20131 16989
rect 20073 16980 20085 16983
rect 19300 16952 20085 16980
rect 19300 16940 19306 16952
rect 20073 16949 20085 16952
rect 20119 16949 20131 16983
rect 20073 16943 20131 16949
rect 552 16890 23368 16912
rect 552 16838 4322 16890
rect 4374 16838 4386 16890
rect 4438 16838 4450 16890
rect 4502 16838 4514 16890
rect 4566 16838 4578 16890
rect 4630 16838 23368 16890
rect 552 16816 23368 16838
rect 4246 16736 4252 16788
rect 4304 16736 4310 16788
rect 5442 16776 5448 16788
rect 4908 16748 5448 16776
rect 4062 16668 4068 16720
rect 4120 16708 4126 16720
rect 4706 16708 4712 16720
rect 4120 16680 4712 16708
rect 4120 16668 4126 16680
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 4908 16717 4936 16748
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 9030 16736 9036 16788
rect 9088 16736 9094 16788
rect 9490 16736 9496 16788
rect 9548 16776 9554 16788
rect 9601 16779 9659 16785
rect 9601 16776 9613 16779
rect 9548 16748 9613 16776
rect 9548 16736 9554 16748
rect 9601 16745 9613 16748
rect 9647 16745 9659 16779
rect 13538 16776 13544 16788
rect 9601 16739 9659 16745
rect 13096 16748 13544 16776
rect 4867 16711 4936 16717
rect 4867 16677 4879 16711
rect 4913 16680 4936 16711
rect 4985 16711 5043 16717
rect 4913 16677 4925 16680
rect 4867 16671 4925 16677
rect 4985 16677 4997 16711
rect 5031 16708 5043 16711
rect 5537 16711 5595 16717
rect 5537 16708 5549 16711
rect 5031 16680 5549 16708
rect 5031 16677 5043 16680
rect 4985 16671 5043 16677
rect 5537 16677 5549 16680
rect 5583 16677 5595 16711
rect 5537 16671 5595 16677
rect 7576 16680 9168 16708
rect 4154 16600 4160 16652
rect 4212 16600 4218 16652
rect 4724 16640 4752 16668
rect 7576 16652 7604 16680
rect 5077 16643 5135 16649
rect 5077 16640 5089 16643
rect 4724 16612 5089 16640
rect 5077 16609 5089 16612
rect 5123 16609 5135 16643
rect 5077 16603 5135 16609
rect 5166 16600 5172 16652
rect 5224 16600 5230 16652
rect 5445 16643 5503 16649
rect 5445 16609 5457 16643
rect 5491 16609 5503 16643
rect 5445 16603 5503 16609
rect 4246 16532 4252 16584
rect 4304 16572 4310 16584
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4304 16544 4629 16572
rect 4304 16532 4310 16544
rect 4617 16541 4629 16544
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 4706 16532 4712 16584
rect 4764 16532 4770 16584
rect 5460 16572 5488 16603
rect 6270 16600 6276 16652
rect 6328 16640 6334 16652
rect 7469 16643 7527 16649
rect 6328 16612 7420 16640
rect 6328 16600 6334 16612
rect 7392 16581 7420 16612
rect 7469 16609 7481 16643
rect 7515 16640 7527 16643
rect 7558 16640 7564 16652
rect 7515 16612 7564 16640
rect 7515 16609 7527 16612
rect 7469 16603 7527 16609
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 8846 16600 8852 16652
rect 8904 16600 8910 16652
rect 9140 16649 9168 16680
rect 9398 16668 9404 16720
rect 9456 16668 9462 16720
rect 9125 16643 9183 16649
rect 9125 16609 9137 16643
rect 9171 16609 9183 16643
rect 9125 16603 9183 16609
rect 9214 16600 9220 16652
rect 9272 16640 9278 16652
rect 13096 16649 13124 16748
rect 13538 16736 13544 16748
rect 13596 16736 13602 16788
rect 14550 16736 14556 16788
rect 14608 16736 14614 16788
rect 15654 16736 15660 16788
rect 15712 16776 15718 16788
rect 16485 16779 16543 16785
rect 15712 16748 16160 16776
rect 15712 16736 15718 16748
rect 13173 16711 13231 16717
rect 13173 16677 13185 16711
rect 13219 16708 13231 16711
rect 14093 16711 14151 16717
rect 13219 16680 13676 16708
rect 13219 16677 13231 16680
rect 13173 16671 13231 16677
rect 9309 16643 9367 16649
rect 9309 16640 9321 16643
rect 9272 16612 9321 16640
rect 9272 16600 9278 16612
rect 9309 16609 9321 16612
rect 9355 16609 9367 16643
rect 9309 16603 9367 16609
rect 13081 16643 13139 16649
rect 13081 16609 13093 16643
rect 13127 16609 13139 16643
rect 13081 16603 13139 16609
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16640 13323 16643
rect 13354 16640 13360 16652
rect 13311 16612 13360 16640
rect 13311 16609 13323 16612
rect 13265 16603 13323 16609
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 13538 16600 13544 16652
rect 13596 16600 13602 16652
rect 13648 16649 13676 16680
rect 14093 16677 14105 16711
rect 14139 16708 14151 16711
rect 14182 16708 14188 16720
rect 14139 16680 14188 16708
rect 14139 16677 14151 16680
rect 14093 16671 14151 16677
rect 14182 16668 14188 16680
rect 14240 16708 14246 16720
rect 14737 16711 14795 16717
rect 14737 16708 14749 16711
rect 14240 16680 14749 16708
rect 14240 16668 14246 16680
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16609 13691 16643
rect 13633 16603 13691 16609
rect 13722 16600 13728 16652
rect 13780 16600 13786 16652
rect 13909 16643 13967 16649
rect 13909 16609 13921 16643
rect 13955 16609 13967 16643
rect 13909 16603 13967 16609
rect 5092 16544 5488 16572
rect 7377 16575 7435 16581
rect 4433 16507 4491 16513
rect 4433 16473 4445 16507
rect 4479 16504 4491 16507
rect 4724 16504 4752 16532
rect 5092 16516 5120 16544
rect 7377 16541 7389 16575
rect 7423 16541 7435 16575
rect 7377 16535 7435 16541
rect 13449 16575 13507 16581
rect 13449 16541 13461 16575
rect 13495 16572 13507 16575
rect 13924 16572 13952 16603
rect 14274 16600 14280 16652
rect 14332 16600 14338 16652
rect 14384 16649 14412 16680
rect 14737 16677 14749 16680
rect 14783 16677 14795 16711
rect 14737 16671 14795 16677
rect 15105 16711 15163 16717
rect 15105 16677 15117 16711
rect 15151 16708 15163 16711
rect 16022 16708 16028 16720
rect 15151 16680 16028 16708
rect 15151 16677 15163 16680
rect 15105 16671 15163 16677
rect 16022 16668 16028 16680
rect 16080 16668 16086 16720
rect 16132 16717 16160 16748
rect 16485 16745 16497 16779
rect 16531 16776 16543 16779
rect 17126 16776 17132 16788
rect 16531 16748 17132 16776
rect 16531 16745 16543 16748
rect 16485 16739 16543 16745
rect 17126 16736 17132 16748
rect 17184 16736 17190 16788
rect 18506 16736 18512 16788
rect 18564 16776 18570 16788
rect 18877 16779 18935 16785
rect 18877 16776 18889 16779
rect 18564 16748 18889 16776
rect 18564 16736 18570 16748
rect 18877 16745 18889 16748
rect 18923 16745 18935 16779
rect 18877 16739 18935 16745
rect 16117 16711 16175 16717
rect 16117 16677 16129 16711
rect 16163 16677 16175 16711
rect 16117 16671 16175 16677
rect 16333 16711 16391 16717
rect 16333 16677 16345 16711
rect 16379 16708 16391 16711
rect 16666 16708 16672 16720
rect 16379 16680 16672 16708
rect 16379 16677 16391 16680
rect 16333 16671 16391 16677
rect 16666 16668 16672 16680
rect 16724 16668 16730 16720
rect 19702 16708 19708 16720
rect 18800 16680 19708 16708
rect 14369 16643 14427 16649
rect 14369 16609 14381 16643
rect 14415 16609 14427 16643
rect 14369 16603 14427 16609
rect 14458 16600 14464 16652
rect 14516 16640 14522 16652
rect 14645 16643 14703 16649
rect 14645 16640 14657 16643
rect 14516 16612 14657 16640
rect 14516 16600 14522 16612
rect 14645 16609 14657 16612
rect 14691 16609 14703 16643
rect 14645 16603 14703 16609
rect 15010 16600 15016 16652
rect 15068 16600 15074 16652
rect 15194 16600 15200 16652
rect 15252 16600 15258 16652
rect 15378 16600 15384 16652
rect 15436 16640 15442 16652
rect 16577 16643 16635 16649
rect 16577 16640 16589 16643
rect 15436 16612 16589 16640
rect 15436 16600 15442 16612
rect 16577 16609 16589 16612
rect 16623 16609 16635 16643
rect 18690 16640 18696 16652
rect 16577 16603 16635 16609
rect 16684 16612 18696 16640
rect 13495 16544 13952 16572
rect 13495 16541 13507 16544
rect 13449 16535 13507 16541
rect 15102 16532 15108 16584
rect 15160 16572 15166 16584
rect 15289 16575 15347 16581
rect 15289 16572 15301 16575
rect 15160 16544 15301 16572
rect 15160 16532 15166 16544
rect 15289 16541 15301 16544
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16572 15531 16575
rect 15654 16572 15660 16584
rect 15519 16544 15660 16572
rect 15519 16541 15531 16544
rect 15473 16535 15531 16541
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 16390 16532 16396 16584
rect 16448 16572 16454 16584
rect 16684 16572 16712 16612
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 18800 16649 18828 16680
rect 19702 16668 19708 16680
rect 19760 16668 19766 16720
rect 21818 16668 21824 16720
rect 21876 16668 21882 16720
rect 18785 16643 18843 16649
rect 18785 16609 18797 16643
rect 18831 16609 18843 16643
rect 18785 16603 18843 16609
rect 18969 16643 19027 16649
rect 18969 16609 18981 16643
rect 19015 16640 19027 16643
rect 19242 16640 19248 16652
rect 19015 16612 19248 16640
rect 19015 16609 19027 16612
rect 18969 16603 19027 16609
rect 18800 16572 18828 16603
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 21542 16600 21548 16652
rect 21600 16600 21606 16652
rect 16448 16544 16712 16572
rect 18064 16544 18828 16572
rect 21821 16575 21879 16581
rect 16448 16532 16454 16544
rect 18064 16516 18092 16544
rect 21821 16541 21833 16575
rect 21867 16572 21879 16575
rect 22094 16572 22100 16584
rect 21867 16544 22100 16572
rect 21867 16541 21879 16544
rect 21821 16535 21879 16541
rect 22094 16532 22100 16544
rect 22152 16572 22158 16584
rect 22554 16572 22560 16584
rect 22152 16544 22560 16572
rect 22152 16532 22158 16544
rect 22554 16532 22560 16544
rect 22612 16532 22618 16584
rect 4479 16476 4752 16504
rect 4479 16473 4491 16476
rect 4433 16467 4491 16473
rect 5074 16464 5080 16516
rect 5132 16464 5138 16516
rect 7837 16507 7895 16513
rect 7837 16473 7849 16507
rect 7883 16504 7895 16507
rect 10226 16504 10232 16516
rect 7883 16476 10232 16504
rect 7883 16473 7895 16476
rect 7837 16467 7895 16473
rect 10226 16464 10232 16476
rect 10284 16464 10290 16516
rect 14921 16507 14979 16513
rect 14921 16473 14933 16507
rect 14967 16504 14979 16507
rect 15562 16504 15568 16516
rect 14967 16476 15568 16504
rect 14967 16473 14979 16476
rect 14921 16467 14979 16473
rect 15562 16464 15568 16476
rect 15620 16464 15626 16516
rect 16206 16464 16212 16516
rect 16264 16504 16270 16516
rect 18046 16504 18052 16516
rect 16264 16476 18052 16504
rect 16264 16464 16270 16476
rect 18046 16464 18052 16476
rect 18104 16464 18110 16516
rect 5350 16396 5356 16448
rect 5408 16396 5414 16448
rect 9585 16439 9643 16445
rect 9585 16405 9597 16439
rect 9631 16436 9643 16439
rect 9674 16436 9680 16448
rect 9631 16408 9680 16436
rect 9631 16405 9643 16408
rect 9585 16399 9643 16405
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 9766 16396 9772 16448
rect 9824 16396 9830 16448
rect 15378 16396 15384 16448
rect 15436 16396 15442 16448
rect 16298 16396 16304 16448
rect 16356 16396 16362 16448
rect 21634 16396 21640 16448
rect 21692 16396 21698 16448
rect 552 16346 23368 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 23368 16346
rect 552 16272 23368 16294
rect 13357 16235 13415 16241
rect 13357 16201 13369 16235
rect 13403 16232 13415 16235
rect 13722 16232 13728 16244
rect 13403 16204 13728 16232
rect 13403 16201 13415 16204
rect 13357 16195 13415 16201
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 15102 16192 15108 16244
rect 15160 16232 15166 16244
rect 16298 16232 16304 16244
rect 15160 16204 16304 16232
rect 15160 16192 15166 16204
rect 16298 16192 16304 16204
rect 16356 16192 16362 16244
rect 16758 16232 16764 16244
rect 16408 16204 16764 16232
rect 6917 16167 6975 16173
rect 6917 16133 6929 16167
rect 6963 16164 6975 16167
rect 7098 16164 7104 16176
rect 6963 16136 7104 16164
rect 6963 16133 6975 16136
rect 6917 16127 6975 16133
rect 7098 16124 7104 16136
rect 7156 16124 7162 16176
rect 12529 16167 12587 16173
rect 12529 16133 12541 16167
rect 12575 16164 12587 16167
rect 12575 16136 13032 16164
rect 12575 16133 12587 16136
rect 12529 16127 12587 16133
rect 5350 16056 5356 16108
rect 5408 16056 5414 16108
rect 5629 16099 5687 16105
rect 5629 16065 5641 16099
rect 5675 16096 5687 16099
rect 6641 16099 6699 16105
rect 6641 16096 6653 16099
rect 5675 16068 6653 16096
rect 5675 16065 5687 16068
rect 5629 16059 5687 16065
rect 6641 16065 6653 16068
rect 6687 16096 6699 16099
rect 6730 16096 6736 16108
rect 6687 16068 6736 16096
rect 6687 16065 6699 16068
rect 6641 16059 6699 16065
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16096 6883 16099
rect 11241 16099 11299 16105
rect 11241 16096 11253 16099
rect 6871 16068 11253 16096
rect 6871 16065 6883 16068
rect 6825 16059 6883 16065
rect 11241 16065 11253 16068
rect 11287 16065 11299 16099
rect 11241 16059 11299 16065
rect 5258 15988 5264 16040
rect 5316 15988 5322 16040
rect 5368 16028 5396 16056
rect 5721 16031 5779 16037
rect 5721 16028 5733 16031
rect 5368 16000 5733 16028
rect 5721 15997 5733 16000
rect 5767 15997 5779 16031
rect 5721 15991 5779 15997
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 15997 5963 16031
rect 5905 15991 5963 15997
rect 6549 16031 6607 16037
rect 6549 15997 6561 16031
rect 6595 16028 6607 16031
rect 7006 16028 7012 16040
rect 6595 16000 7012 16028
rect 6595 15997 6607 16000
rect 6549 15991 6607 15997
rect 5276 15960 5304 15988
rect 5920 15960 5948 15991
rect 7006 15988 7012 16000
rect 7064 16028 7070 16040
rect 7101 16031 7159 16037
rect 7101 16028 7113 16031
rect 7064 16000 7113 16028
rect 7064 15988 7070 16000
rect 7101 15997 7113 16000
rect 7147 15997 7159 16031
rect 7101 15991 7159 15997
rect 5276 15932 5948 15960
rect 6914 15920 6920 15972
rect 6972 15920 6978 15972
rect 7116 15960 7144 15991
rect 7190 15988 7196 16040
rect 7248 15988 7254 16040
rect 8018 15960 8024 15972
rect 7116 15932 8024 15960
rect 8018 15920 8024 15932
rect 8076 15920 8082 15972
rect 11256 15960 11284 16059
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11664 16068 11713 16096
rect 11664 16056 11670 16068
rect 11701 16065 11713 16068
rect 11747 16096 11759 16099
rect 11747 16068 12296 16096
rect 11747 16065 11759 16068
rect 11701 16059 11759 16065
rect 11333 16031 11391 16037
rect 11333 15997 11345 16031
rect 11379 16028 11391 16031
rect 11422 16028 11428 16040
rect 11379 16000 11428 16028
rect 11379 15997 11391 16000
rect 11333 15991 11391 15997
rect 11422 15988 11428 16000
rect 11480 16028 11486 16040
rect 12268 16037 12296 16068
rect 11793 16031 11851 16037
rect 11793 16028 11805 16031
rect 11480 16000 11805 16028
rect 11480 15988 11486 16000
rect 11793 15997 11805 16000
rect 11839 15997 11851 16031
rect 11793 15991 11851 15997
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 15997 12311 16031
rect 12253 15991 12311 15997
rect 11992 15960 12020 15991
rect 13004 15972 13032 16136
rect 13538 16124 13544 16176
rect 13596 16164 13602 16176
rect 14461 16167 14519 16173
rect 13596 16136 13676 16164
rect 13596 16124 13602 16136
rect 13354 16056 13360 16108
rect 13412 16096 13418 16108
rect 13648 16105 13676 16136
rect 14461 16133 14473 16167
rect 14507 16164 14519 16167
rect 15194 16164 15200 16176
rect 14507 16136 15200 16164
rect 14507 16133 14519 16136
rect 14461 16127 14519 16133
rect 15194 16124 15200 16136
rect 15252 16164 15258 16176
rect 15381 16167 15439 16173
rect 15381 16164 15393 16167
rect 15252 16136 15393 16164
rect 15252 16124 15258 16136
rect 15381 16133 15393 16136
rect 15427 16133 15439 16167
rect 16408 16164 16436 16204
rect 16758 16192 16764 16204
rect 16816 16192 16822 16244
rect 18598 16192 18604 16244
rect 18656 16232 18662 16244
rect 19153 16235 19211 16241
rect 19153 16232 19165 16235
rect 18656 16204 19165 16232
rect 18656 16192 18662 16204
rect 19153 16201 19165 16204
rect 19199 16232 19211 16235
rect 19426 16232 19432 16244
rect 19199 16204 19432 16232
rect 19199 16201 19211 16204
rect 19153 16195 19211 16201
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 21542 16192 21548 16244
rect 21600 16192 21606 16244
rect 21821 16235 21879 16241
rect 21821 16201 21833 16235
rect 21867 16232 21879 16235
rect 22094 16232 22100 16244
rect 21867 16204 22100 16232
rect 21867 16201 21879 16204
rect 21821 16195 21879 16201
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 22557 16235 22615 16241
rect 22557 16201 22569 16235
rect 22603 16232 22615 16235
rect 22646 16232 22652 16244
rect 22603 16204 22652 16232
rect 22603 16201 22615 16204
rect 22557 16195 22615 16201
rect 22646 16192 22652 16204
rect 22704 16192 22710 16244
rect 15381 16127 15439 16133
rect 16132 16136 16436 16164
rect 13633 16099 13691 16105
rect 13412 16068 13584 16096
rect 13412 16056 13418 16068
rect 13173 16031 13231 16037
rect 13173 15997 13185 16031
rect 13219 16028 13231 16031
rect 13446 16028 13452 16040
rect 13219 16000 13452 16028
rect 13219 15997 13231 16000
rect 13173 15991 13231 15997
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 13556 16028 13584 16068
rect 13633 16065 13645 16099
rect 13679 16065 13691 16099
rect 13633 16059 13691 16065
rect 15102 16056 15108 16108
rect 15160 16096 15166 16108
rect 15289 16099 15347 16105
rect 15289 16096 15301 16099
rect 15160 16068 15301 16096
rect 15160 16056 15166 16068
rect 15289 16065 15301 16068
rect 15335 16065 15347 16099
rect 15654 16096 15660 16108
rect 15289 16059 15347 16065
rect 15488 16068 15660 16096
rect 13725 16031 13783 16037
rect 13725 16028 13737 16031
rect 13556 16000 13737 16028
rect 13725 15997 13737 16000
rect 13771 15997 13783 16031
rect 13725 15991 13783 15997
rect 14182 15988 14188 16040
rect 14240 15988 14246 16040
rect 14461 16031 14519 16037
rect 14461 15997 14473 16031
rect 14507 16028 14519 16031
rect 15010 16028 15016 16040
rect 14507 16000 15016 16028
rect 14507 15997 14519 16000
rect 14461 15991 14519 15997
rect 15010 15988 15016 16000
rect 15068 15988 15074 16040
rect 15194 15988 15200 16040
rect 15252 15988 15258 16040
rect 15488 16037 15516 16068
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 16132 16104 16160 16136
rect 16666 16124 16672 16176
rect 16724 16124 16730 16176
rect 16942 16124 16948 16176
rect 17000 16124 17006 16176
rect 19518 16164 19524 16176
rect 19260 16136 19524 16164
rect 16132 16076 16252 16104
rect 15473 16031 15531 16037
rect 15473 15997 15485 16031
rect 15519 15997 15531 16031
rect 15473 15991 15531 15997
rect 16114 15988 16120 16040
rect 16172 15988 16178 16040
rect 16224 16037 16252 16076
rect 16298 16056 16304 16108
rect 16356 16056 16362 16108
rect 16393 16099 16451 16105
rect 16393 16065 16405 16099
rect 16439 16096 16451 16099
rect 16684 16096 16712 16124
rect 19260 16096 19288 16136
rect 19518 16124 19524 16136
rect 19576 16124 19582 16176
rect 19702 16124 19708 16176
rect 19760 16164 19766 16176
rect 19797 16167 19855 16173
rect 19797 16164 19809 16167
rect 19760 16136 19809 16164
rect 19760 16124 19766 16136
rect 19797 16133 19809 16136
rect 19843 16133 19855 16167
rect 21560 16164 21588 16192
rect 19797 16127 19855 16133
rect 21192 16136 21772 16164
rect 16439 16068 16988 16096
rect 16439 16065 16451 16068
rect 16393 16059 16451 16065
rect 16209 16031 16267 16037
rect 16209 15997 16221 16031
rect 16255 15997 16267 16031
rect 16316 16028 16344 16056
rect 16482 16028 16488 16040
rect 16316 16000 16488 16028
rect 16209 15991 16267 15997
rect 16482 15988 16488 16000
rect 16540 16028 16546 16040
rect 16669 16031 16727 16037
rect 16669 16028 16681 16031
rect 16540 16000 16681 16028
rect 16540 15988 16546 16000
rect 16669 15997 16681 16000
rect 16715 15997 16727 16031
rect 16669 15991 16727 15997
rect 16758 15988 16764 16040
rect 16816 15988 16822 16040
rect 16960 16037 16988 16068
rect 19168 16068 19288 16096
rect 19168 16040 19196 16068
rect 19426 16056 19432 16108
rect 19484 16096 19490 16108
rect 19613 16099 19671 16105
rect 19613 16096 19625 16099
rect 19484 16068 19625 16096
rect 19484 16056 19490 16068
rect 19613 16065 19625 16068
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 19720 16068 19932 16096
rect 16945 16031 17003 16037
rect 16945 15997 16957 16031
rect 16991 15997 17003 16031
rect 16945 15991 17003 15997
rect 19150 15988 19156 16040
rect 19208 15988 19214 16040
rect 19242 15988 19248 16040
rect 19300 16028 19306 16040
rect 19720 16028 19748 16068
rect 19904 16037 19932 16068
rect 20364 16068 20760 16096
rect 20364 16040 20392 16068
rect 19300 16000 19748 16028
rect 19889 16031 19947 16037
rect 19300 15988 19306 16000
rect 19889 15997 19901 16031
rect 19935 15997 19947 16031
rect 19889 15991 19947 15997
rect 20257 16031 20315 16037
rect 20257 15997 20269 16031
rect 20303 16028 20315 16031
rect 20346 16028 20352 16040
rect 20303 16000 20352 16028
rect 20303 15997 20315 16000
rect 20257 15991 20315 15997
rect 20346 15988 20352 16000
rect 20404 15988 20410 16040
rect 20732 16037 20760 16068
rect 21192 16037 21220 16136
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 20717 16031 20775 16037
rect 20717 15997 20729 16031
rect 20763 15997 20775 16031
rect 20717 15991 20775 15997
rect 21177 16031 21235 16037
rect 21177 15997 21189 16031
rect 21223 15997 21235 16031
rect 21177 15991 21235 15997
rect 21284 16028 21312 16059
rect 21450 16056 21456 16108
rect 21508 16096 21514 16108
rect 21744 16105 21772 16136
rect 21545 16099 21603 16105
rect 21545 16096 21557 16099
rect 21508 16068 21557 16096
rect 21508 16056 21514 16068
rect 21545 16065 21557 16068
rect 21591 16065 21603 16099
rect 21545 16059 21603 16065
rect 21729 16099 21787 16105
rect 21729 16065 21741 16099
rect 21775 16065 21787 16099
rect 21729 16059 21787 16065
rect 22186 16056 22192 16108
rect 22244 16056 22250 16108
rect 21634 16028 21640 16040
rect 21284 16000 21640 16028
rect 11256 15932 12020 15960
rect 12161 15963 12219 15969
rect 12161 15929 12173 15963
rect 12207 15960 12219 15963
rect 12529 15963 12587 15969
rect 12529 15960 12541 15963
rect 12207 15932 12541 15960
rect 12207 15929 12219 15932
rect 12161 15923 12219 15929
rect 12529 15929 12541 15932
rect 12575 15929 12587 15963
rect 12529 15923 12587 15929
rect 12986 15920 12992 15972
rect 13044 15920 13050 15972
rect 15657 15963 15715 15969
rect 15657 15929 15669 15963
rect 15703 15960 15715 15963
rect 20073 15963 20131 15969
rect 20073 15960 20085 15963
rect 15703 15932 16712 15960
rect 15703 15929 15715 15932
rect 15657 15923 15715 15929
rect 16684 15904 16712 15932
rect 19536 15932 20085 15960
rect 19536 15904 19564 15932
rect 20073 15929 20085 15932
rect 20119 15960 20131 15963
rect 20548 15960 20576 15991
rect 20806 15960 20812 15972
rect 20119 15932 20576 15960
rect 20640 15932 20812 15960
rect 20119 15929 20131 15932
rect 20073 15923 20131 15929
rect 5905 15895 5963 15901
rect 5905 15861 5917 15895
rect 5951 15892 5963 15895
rect 6181 15895 6239 15901
rect 6181 15892 6193 15895
rect 5951 15864 6193 15892
rect 5951 15861 5963 15864
rect 5905 15855 5963 15861
rect 6181 15861 6193 15864
rect 6227 15861 6239 15895
rect 6181 15855 6239 15861
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 11698 15892 11704 15904
rect 11480 15864 11704 15892
rect 11480 15852 11486 15864
rect 11698 15852 11704 15864
rect 11756 15892 11762 15904
rect 12345 15895 12403 15901
rect 12345 15892 12357 15895
rect 11756 15864 12357 15892
rect 11756 15852 11762 15864
rect 12345 15861 12357 15864
rect 12391 15861 12403 15895
rect 12345 15855 12403 15861
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 14093 15895 14151 15901
rect 14093 15892 14105 15895
rect 13596 15864 14105 15892
rect 13596 15852 13602 15864
rect 14093 15861 14105 15864
rect 14139 15861 14151 15895
rect 14093 15855 14151 15861
rect 14274 15852 14280 15904
rect 14332 15852 14338 15904
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 16298 15892 16304 15904
rect 15436 15864 16304 15892
rect 15436 15852 15442 15864
rect 16298 15852 16304 15864
rect 16356 15852 16362 15904
rect 16574 15852 16580 15904
rect 16632 15852 16638 15904
rect 16666 15852 16672 15904
rect 16724 15852 16730 15904
rect 19518 15852 19524 15904
rect 19576 15852 19582 15904
rect 19613 15895 19671 15901
rect 19613 15861 19625 15895
rect 19659 15892 19671 15895
rect 19702 15892 19708 15904
rect 19659 15864 19708 15892
rect 19659 15861 19671 15864
rect 19613 15855 19671 15861
rect 19702 15852 19708 15864
rect 19760 15852 19766 15904
rect 20441 15895 20499 15901
rect 20441 15861 20453 15895
rect 20487 15892 20499 15895
rect 20640 15892 20668 15932
rect 20806 15920 20812 15932
rect 20864 15960 20870 15972
rect 21284 15960 21312 16000
rect 21634 15988 21640 16000
rect 21692 15988 21698 16040
rect 22204 16028 22232 16056
rect 22373 16031 22431 16037
rect 22373 16028 22385 16031
rect 22204 16000 22385 16028
rect 22373 15997 22385 16000
rect 22419 15997 22431 16031
rect 22373 15991 22431 15997
rect 20864 15932 21312 15960
rect 22189 15963 22247 15969
rect 20864 15920 20870 15932
rect 22189 15929 22201 15963
rect 22235 15929 22247 15963
rect 22189 15923 22247 15929
rect 20487 15864 20668 15892
rect 20487 15861 20499 15864
rect 20441 15855 20499 15861
rect 20714 15852 20720 15904
rect 20772 15852 20778 15904
rect 21634 15852 21640 15904
rect 21692 15892 21698 15904
rect 22005 15895 22063 15901
rect 22005 15892 22017 15895
rect 21692 15864 22017 15892
rect 21692 15852 21698 15864
rect 22005 15861 22017 15864
rect 22051 15892 22063 15895
rect 22204 15892 22232 15923
rect 22051 15864 22232 15892
rect 22051 15861 22063 15864
rect 22005 15855 22063 15861
rect 552 15802 23368 15824
rect 552 15750 4322 15802
rect 4374 15750 4386 15802
rect 4438 15750 4450 15802
rect 4502 15750 4514 15802
rect 4566 15750 4578 15802
rect 4630 15750 23368 15802
rect 552 15728 23368 15750
rect 4246 15648 4252 15700
rect 4304 15688 4310 15700
rect 4433 15691 4491 15697
rect 4433 15688 4445 15691
rect 4304 15660 4445 15688
rect 4304 15648 4310 15660
rect 4433 15657 4445 15660
rect 4479 15688 4491 15691
rect 4798 15688 4804 15700
rect 4479 15660 4804 15688
rect 4479 15657 4491 15660
rect 4433 15651 4491 15657
rect 4798 15648 4804 15660
rect 4856 15648 4862 15700
rect 15194 15648 15200 15700
rect 15252 15688 15258 15700
rect 20162 15688 20168 15700
rect 15252 15660 20168 15688
rect 15252 15648 15258 15660
rect 20162 15648 20168 15660
rect 20220 15648 20226 15700
rect 20806 15648 20812 15700
rect 20864 15648 20870 15700
rect 10134 15620 10140 15632
rect 8772 15592 9352 15620
rect 4062 15512 4068 15564
rect 4120 15512 4126 15564
rect 4249 15555 4307 15561
rect 4249 15521 4261 15555
rect 4295 15552 4307 15555
rect 5074 15552 5080 15564
rect 4295 15524 5080 15552
rect 4295 15521 4307 15524
rect 4249 15515 4307 15521
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 5261 15555 5319 15561
rect 5261 15521 5273 15555
rect 5307 15552 5319 15555
rect 5810 15552 5816 15564
rect 5307 15524 5816 15552
rect 5307 15521 5319 15524
rect 5261 15515 5319 15521
rect 5810 15512 5816 15524
rect 5868 15512 5874 15564
rect 5994 15512 6000 15564
rect 6052 15512 6058 15564
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15552 6699 15555
rect 7285 15555 7343 15561
rect 7285 15552 7297 15555
rect 6687 15524 7297 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 7285 15521 7297 15524
rect 7331 15552 7343 15555
rect 7558 15552 7564 15564
rect 7331 15524 7564 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 7558 15512 7564 15524
rect 7616 15512 7622 15564
rect 4706 15444 4712 15496
rect 4764 15484 4770 15496
rect 5169 15487 5227 15493
rect 5169 15484 5181 15487
rect 4764 15456 5181 15484
rect 4764 15444 4770 15456
rect 5169 15453 5181 15456
rect 5215 15453 5227 15487
rect 5169 15447 5227 15453
rect 6086 15444 6092 15496
rect 6144 15444 6150 15496
rect 6730 15444 6736 15496
rect 6788 15444 6794 15496
rect 7190 15484 7196 15496
rect 6932 15456 7196 15484
rect 5629 15419 5687 15425
rect 5629 15385 5641 15419
rect 5675 15416 5687 15419
rect 5994 15416 6000 15428
rect 5675 15388 6000 15416
rect 5675 15385 5687 15388
rect 5629 15379 5687 15385
rect 5994 15376 6000 15388
rect 6052 15376 6058 15428
rect 6365 15419 6423 15425
rect 6365 15385 6377 15419
rect 6411 15416 6423 15419
rect 6932 15416 6960 15456
rect 7190 15444 7196 15456
rect 7248 15444 7254 15496
rect 8662 15444 8668 15496
rect 8720 15484 8726 15496
rect 8772 15493 8800 15592
rect 9324 15561 9352 15592
rect 9968 15592 10140 15620
rect 9968 15561 9996 15592
rect 10134 15580 10140 15592
rect 10192 15620 10198 15632
rect 11514 15620 11520 15632
rect 10192 15592 11520 15620
rect 10192 15580 10198 15592
rect 11514 15580 11520 15592
rect 11572 15580 11578 15632
rect 16482 15580 16488 15632
rect 16540 15580 16546 15632
rect 16574 15580 16580 15632
rect 16632 15620 16638 15632
rect 20257 15623 20315 15629
rect 16632 15592 17080 15620
rect 16632 15580 16638 15592
rect 8849 15555 8907 15561
rect 8849 15521 8861 15555
rect 8895 15521 8907 15555
rect 8849 15515 8907 15521
rect 9309 15555 9367 15561
rect 9309 15521 9321 15555
rect 9355 15521 9367 15555
rect 9309 15515 9367 15521
rect 9402 15555 9460 15561
rect 9402 15521 9414 15555
rect 9448 15521 9460 15555
rect 9402 15515 9460 15521
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15521 10011 15555
rect 9953 15515 10011 15521
rect 10046 15555 10104 15561
rect 10046 15521 10058 15555
rect 10092 15521 10104 15555
rect 10046 15515 10104 15521
rect 8757 15487 8815 15493
rect 8757 15484 8769 15487
rect 8720 15456 8769 15484
rect 8720 15444 8726 15456
rect 8757 15453 8769 15456
rect 8803 15453 8815 15487
rect 8757 15447 8815 15453
rect 8864 15484 8892 15515
rect 9416 15484 9444 15515
rect 10060 15484 10088 15515
rect 11422 15512 11428 15564
rect 11480 15552 11486 15564
rect 11701 15555 11759 15561
rect 11701 15552 11713 15555
rect 11480 15524 11713 15552
rect 11480 15512 11486 15524
rect 11701 15521 11713 15524
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 12986 15512 12992 15564
rect 13044 15512 13050 15564
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 13446 15552 13452 15564
rect 13403 15524 13452 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 13446 15512 13452 15524
rect 13504 15512 13510 15564
rect 16206 15512 16212 15564
rect 16264 15552 16270 15564
rect 16301 15555 16359 15561
rect 16301 15552 16313 15555
rect 16264 15524 16313 15552
rect 16264 15512 16270 15524
rect 16301 15521 16313 15524
rect 16347 15521 16359 15555
rect 16301 15515 16359 15521
rect 16393 15555 16451 15561
rect 16393 15521 16405 15555
rect 16439 15521 16451 15555
rect 16393 15515 16451 15521
rect 8864 15456 9444 15484
rect 9692 15456 10088 15484
rect 6411 15388 6960 15416
rect 6411 15385 6423 15388
rect 6365 15379 6423 15385
rect 7006 15376 7012 15428
rect 7064 15376 7070 15428
rect 7653 15419 7711 15425
rect 7653 15385 7665 15419
rect 7699 15416 7711 15419
rect 8864 15416 8892 15456
rect 9692 15428 9720 15456
rect 11606 15444 11612 15496
rect 11664 15444 11670 15496
rect 13814 15444 13820 15496
rect 13872 15484 13878 15496
rect 13909 15487 13967 15493
rect 13909 15484 13921 15487
rect 13872 15456 13921 15484
rect 13872 15444 13878 15456
rect 13909 15453 13921 15456
rect 13955 15453 13967 15487
rect 16408 15484 16436 15515
rect 16666 15512 16672 15564
rect 16724 15512 16730 15564
rect 16942 15512 16948 15564
rect 17000 15512 17006 15564
rect 17052 15561 17080 15592
rect 20257 15589 20269 15623
rect 20303 15589 20315 15623
rect 20257 15583 20315 15589
rect 20473 15623 20531 15629
rect 20473 15589 20485 15623
rect 20519 15620 20531 15623
rect 20519 15592 20760 15620
rect 20519 15589 20531 15592
rect 20473 15583 20531 15589
rect 17037 15555 17095 15561
rect 17037 15521 17049 15555
rect 17083 15521 17095 15555
rect 17037 15515 17095 15521
rect 17310 15512 17316 15564
rect 17368 15512 17374 15564
rect 19518 15512 19524 15564
rect 19576 15512 19582 15564
rect 19702 15512 19708 15564
rect 19760 15512 19766 15564
rect 16850 15484 16856 15496
rect 16408 15456 16856 15484
rect 13909 15447 13967 15453
rect 16850 15444 16856 15456
rect 16908 15444 16914 15496
rect 20272 15484 20300 15583
rect 20732 15564 20760 15592
rect 20714 15512 20720 15564
rect 20772 15512 20778 15564
rect 20993 15555 21051 15561
rect 20993 15521 21005 15555
rect 21039 15521 21051 15555
rect 20993 15515 21051 15521
rect 21729 15555 21787 15561
rect 21729 15521 21741 15555
rect 21775 15552 21787 15555
rect 22186 15552 22192 15564
rect 21775 15524 22192 15552
rect 21775 15521 21787 15524
rect 21729 15515 21787 15521
rect 21008 15484 21036 15515
rect 22186 15512 22192 15524
rect 22244 15512 22250 15564
rect 20272 15456 21036 15484
rect 7699 15388 8892 15416
rect 9217 15419 9275 15425
rect 7699 15385 7711 15388
rect 7653 15379 7711 15385
rect 9217 15385 9229 15419
rect 9263 15416 9275 15419
rect 9674 15416 9680 15428
rect 9263 15388 9680 15416
rect 9263 15385 9275 15388
rect 9217 15379 9275 15385
rect 9674 15376 9680 15388
rect 9732 15376 9738 15428
rect 12066 15376 12072 15428
rect 12124 15376 12130 15428
rect 20806 15416 20812 15428
rect 20456 15388 20812 15416
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 9950 15348 9956 15360
rect 9539 15320 9956 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 9950 15308 9956 15320
rect 10008 15308 10014 15360
rect 10042 15308 10048 15360
rect 10100 15348 10106 15360
rect 10137 15351 10195 15357
rect 10137 15348 10149 15351
rect 10100 15320 10149 15348
rect 10100 15308 10106 15320
rect 10137 15317 10149 15320
rect 10183 15317 10195 15351
rect 10137 15311 10195 15317
rect 15930 15308 15936 15360
rect 15988 15348 15994 15360
rect 16117 15351 16175 15357
rect 16117 15348 16129 15351
rect 15988 15320 16129 15348
rect 15988 15308 15994 15320
rect 16117 15317 16129 15320
rect 16163 15317 16175 15351
rect 16117 15311 16175 15317
rect 16758 15308 16764 15360
rect 16816 15308 16822 15360
rect 17126 15308 17132 15360
rect 17184 15348 17190 15360
rect 17221 15351 17279 15357
rect 17221 15348 17233 15351
rect 17184 15320 17233 15348
rect 17184 15308 17190 15320
rect 17221 15317 17233 15320
rect 17267 15348 17279 15351
rect 18782 15348 18788 15360
rect 17267 15320 18788 15348
rect 17267 15317 17279 15320
rect 17221 15311 17279 15317
rect 18782 15308 18788 15320
rect 18840 15308 18846 15360
rect 19613 15351 19671 15357
rect 19613 15317 19625 15351
rect 19659 15348 19671 15351
rect 19702 15348 19708 15360
rect 19659 15320 19708 15348
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 20456 15357 20484 15388
rect 20806 15376 20812 15388
rect 20864 15376 20870 15428
rect 20441 15351 20499 15357
rect 20441 15317 20453 15351
rect 20487 15317 20499 15351
rect 20441 15311 20499 15317
rect 20530 15308 20536 15360
rect 20588 15348 20594 15360
rect 20625 15351 20683 15357
rect 20625 15348 20637 15351
rect 20588 15320 20637 15348
rect 20588 15308 20594 15320
rect 20625 15317 20637 15320
rect 20671 15317 20683 15351
rect 20625 15311 20683 15317
rect 20714 15308 20720 15360
rect 20772 15348 20778 15360
rect 20916 15348 20944 15456
rect 21634 15444 21640 15496
rect 21692 15444 21698 15496
rect 20772 15320 20944 15348
rect 20772 15308 20778 15320
rect 20990 15308 20996 15360
rect 21048 15308 21054 15360
rect 22094 15308 22100 15360
rect 22152 15308 22158 15360
rect 552 15258 23368 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 23368 15258
rect 552 15184 23368 15206
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 6549 15147 6607 15153
rect 4212 15116 5396 15144
rect 4212 15104 4218 15116
rect 5077 15079 5135 15085
rect 5077 15045 5089 15079
rect 5123 15045 5135 15079
rect 5077 15039 5135 15045
rect 4632 14980 4936 15008
rect 4632 14949 4660 14980
rect 4617 14943 4675 14949
rect 4617 14909 4629 14943
rect 4663 14909 4675 14943
rect 4617 14903 4675 14909
rect 4798 14900 4804 14952
rect 4856 14900 4862 14952
rect 4709 14875 4767 14881
rect 4709 14841 4721 14875
rect 4755 14841 4767 14875
rect 4908 14872 4936 14980
rect 4985 14943 5043 14949
rect 4985 14909 4997 14943
rect 5031 14940 5043 14943
rect 5092 14940 5120 15039
rect 5031 14912 5120 14940
rect 5031 14909 5043 14912
rect 4985 14903 5043 14909
rect 5166 14900 5172 14952
rect 5224 14940 5230 14952
rect 5368 14949 5396 15116
rect 6549 15113 6561 15147
rect 6595 15144 6607 15147
rect 6914 15144 6920 15156
rect 6595 15116 6920 15144
rect 6595 15113 6607 15116
rect 6549 15107 6607 15113
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 7190 15104 7196 15156
rect 7248 15144 7254 15156
rect 11882 15144 11888 15156
rect 7248 15116 11888 15144
rect 7248 15104 7254 15116
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 12713 15147 12771 15153
rect 12713 15144 12725 15147
rect 12406 15116 12725 15144
rect 5994 15036 6000 15088
rect 6052 15076 6058 15088
rect 6365 15079 6423 15085
rect 6365 15076 6377 15079
rect 6052 15048 6377 15076
rect 6052 15036 6058 15048
rect 6365 15045 6377 15048
rect 6411 15045 6423 15079
rect 6365 15039 6423 15045
rect 7929 15079 7987 15085
rect 7929 15045 7941 15079
rect 7975 15076 7987 15079
rect 7975 15048 10548 15076
rect 7975 15045 7987 15048
rect 7929 15039 7987 15045
rect 6086 14968 6092 15020
rect 6144 14968 6150 15020
rect 7098 15008 7104 15020
rect 6932 14980 7104 15008
rect 5261 14943 5319 14949
rect 5261 14940 5273 14943
rect 5224 14912 5273 14940
rect 5224 14900 5230 14912
rect 5261 14909 5273 14912
rect 5307 14909 5319 14943
rect 5261 14903 5319 14909
rect 5353 14943 5411 14949
rect 5353 14909 5365 14943
rect 5399 14940 5411 14943
rect 5442 14940 5448 14952
rect 5399 14912 5448 14940
rect 5399 14909 5411 14912
rect 5353 14903 5411 14909
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 6932 14949 6960 14980
rect 7098 14968 7104 14980
rect 7156 15008 7162 15020
rect 7469 15011 7527 15017
rect 7469 15008 7481 15011
rect 7156 14980 7481 15008
rect 7156 14968 7162 14980
rect 7469 14977 7481 14980
rect 7515 14977 7527 15011
rect 7469 14971 7527 14977
rect 9674 14968 9680 15020
rect 9732 14968 9738 15020
rect 10520 15017 10548 15048
rect 10505 15011 10563 15017
rect 10505 14977 10517 15011
rect 10551 15008 10563 15011
rect 11425 15011 11483 15017
rect 10551 14980 11376 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14909 6975 14943
rect 6917 14903 6975 14909
rect 7006 14900 7012 14952
rect 7064 14940 7070 14952
rect 7561 14943 7619 14949
rect 7561 14940 7573 14943
rect 7064 14912 7573 14940
rect 7064 14900 7070 14912
rect 7561 14909 7573 14912
rect 7607 14909 7619 14943
rect 7561 14903 7619 14909
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14940 9827 14943
rect 10134 14940 10140 14952
rect 9815 14912 10140 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 10134 14900 10140 14912
rect 10192 14900 10198 14952
rect 10597 14943 10655 14949
rect 10597 14909 10609 14943
rect 10643 14940 10655 14943
rect 11238 14940 11244 14952
rect 10643 14912 11244 14940
rect 10643 14909 10655 14912
rect 10597 14903 10655 14909
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 11348 14949 11376 14980
rect 11425 14977 11437 15011
rect 11471 15008 11483 15011
rect 12406 15008 12434 15116
rect 12713 15113 12725 15116
rect 12759 15113 12771 15147
rect 12713 15107 12771 15113
rect 14093 15147 14151 15153
rect 14093 15113 14105 15147
rect 14139 15144 14151 15147
rect 14274 15144 14280 15156
rect 14139 15116 14280 15144
rect 14139 15113 14151 15116
rect 14093 15107 14151 15113
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 14384 15116 16620 15144
rect 12802 15036 12808 15088
rect 12860 15076 12866 15088
rect 14384 15076 14412 15116
rect 12860 15048 14412 15076
rect 16592 15076 16620 15116
rect 16850 15104 16856 15156
rect 16908 15144 16914 15156
rect 17034 15144 17040 15156
rect 16908 15116 17040 15144
rect 16908 15104 16914 15116
rect 17034 15104 17040 15116
rect 17092 15104 17098 15156
rect 18233 15147 18291 15153
rect 18233 15113 18245 15147
rect 18279 15144 18291 15147
rect 18690 15144 18696 15156
rect 18279 15116 18696 15144
rect 18279 15113 18291 15116
rect 18233 15107 18291 15113
rect 18690 15104 18696 15116
rect 18748 15104 18754 15156
rect 20533 15147 20591 15153
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 20990 15144 20996 15156
rect 20579 15116 20996 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 20717 15079 20775 15085
rect 16592 15048 20668 15076
rect 12860 15036 12866 15048
rect 11471 14980 12434 15008
rect 17865 15011 17923 15017
rect 11471 14977 11483 14980
rect 11425 14971 11483 14977
rect 11333 14943 11391 14949
rect 11333 14909 11345 14943
rect 11379 14909 11391 14943
rect 11333 14903 11391 14909
rect 11514 14900 11520 14952
rect 11572 14900 11578 14952
rect 11992 14949 12020 14980
rect 17865 14977 17877 15011
rect 17911 15008 17923 15011
rect 17911 14980 18092 15008
rect 17911 14977 17923 14980
rect 17865 14971 17923 14977
rect 18064 14952 18092 14980
rect 18598 14968 18604 15020
rect 18656 15008 18662 15020
rect 18693 15011 18751 15017
rect 18693 15008 18705 15011
rect 18656 14980 18705 15008
rect 18656 14968 18662 14980
rect 18693 14977 18705 14980
rect 18739 14977 18751 15011
rect 19150 15008 19156 15020
rect 18693 14971 18751 14977
rect 18800 14980 19156 15008
rect 11977 14943 12035 14949
rect 11977 14909 11989 14943
rect 12023 14909 12035 14943
rect 11977 14903 12035 14909
rect 12066 14900 12072 14952
rect 12124 14940 12130 14952
rect 12253 14943 12311 14949
rect 12253 14940 12265 14943
rect 12124 14912 12265 14940
rect 12124 14900 12130 14912
rect 12253 14909 12265 14912
rect 12299 14940 12311 14943
rect 12299 14912 12664 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 5077 14875 5135 14881
rect 5077 14872 5089 14875
rect 4908 14844 5089 14872
rect 4709 14835 4767 14841
rect 5077 14841 5089 14844
rect 5123 14872 5135 14875
rect 7285 14875 7343 14881
rect 5123 14844 6960 14872
rect 5123 14841 5135 14844
rect 5077 14835 5135 14841
rect 4246 14764 4252 14816
rect 4304 14804 4310 14816
rect 4433 14807 4491 14813
rect 4433 14804 4445 14807
rect 4304 14776 4445 14804
rect 4304 14764 4310 14776
rect 4433 14773 4445 14776
rect 4479 14773 4491 14807
rect 4724 14804 4752 14835
rect 6932 14816 6960 14844
rect 7285 14841 7297 14875
rect 7331 14872 7343 14875
rect 12529 14875 12587 14881
rect 12529 14872 12541 14875
rect 7331 14844 12541 14872
rect 7331 14841 7343 14844
rect 7285 14835 7343 14841
rect 5626 14804 5632 14816
rect 4724 14776 5632 14804
rect 4433 14767 4491 14773
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 6914 14764 6920 14816
rect 6972 14764 6978 14816
rect 9401 14807 9459 14813
rect 9401 14773 9413 14807
rect 9447 14804 9459 14807
rect 9674 14804 9680 14816
rect 9447 14776 9680 14804
rect 9447 14773 9459 14776
rect 9401 14767 9459 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 10229 14807 10287 14813
rect 10229 14773 10241 14807
rect 10275 14804 10287 14807
rect 10318 14804 10324 14816
rect 10275 14776 10324 14804
rect 10275 14773 10287 14776
rect 10229 14767 10287 14773
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 12084 14813 12112 14844
rect 12529 14841 12541 14844
rect 12575 14841 12587 14875
rect 12636 14872 12664 14912
rect 13538 14900 13544 14952
rect 13596 14900 13602 14952
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13722 14940 13728 14952
rect 13679 14912 13728 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 15930 14949 15936 14952
rect 13817 14943 13875 14949
rect 13817 14909 13829 14943
rect 13863 14909 13875 14943
rect 13817 14903 13875 14909
rect 13909 14943 13967 14949
rect 13909 14909 13921 14943
rect 13955 14909 13967 14943
rect 13909 14903 13967 14909
rect 15657 14943 15715 14949
rect 15657 14909 15669 14943
rect 15703 14909 15715 14943
rect 15924 14940 15936 14949
rect 15891 14912 15936 14940
rect 15657 14903 15715 14909
rect 15924 14903 15936 14912
rect 12729 14875 12787 14881
rect 12729 14872 12741 14875
rect 12636 14844 12741 14872
rect 12529 14835 12587 14841
rect 12729 14841 12741 14844
rect 12775 14841 12787 14875
rect 13832 14872 13860 14903
rect 12729 14835 12787 14841
rect 12820 14844 13860 14872
rect 12069 14807 12127 14813
rect 12069 14773 12081 14807
rect 12115 14773 12127 14807
rect 12069 14767 12127 14773
rect 12158 14764 12164 14816
rect 12216 14804 12222 14816
rect 12437 14807 12495 14813
rect 12437 14804 12449 14807
rect 12216 14776 12449 14804
rect 12216 14764 12222 14776
rect 12437 14773 12449 14776
rect 12483 14804 12495 14807
rect 12820 14804 12848 14844
rect 12483 14776 12848 14804
rect 12897 14807 12955 14813
rect 12483 14773 12495 14776
rect 12437 14767 12495 14773
rect 12897 14773 12909 14807
rect 12943 14804 12955 14807
rect 13170 14804 13176 14816
rect 12943 14776 13176 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 13722 14764 13728 14816
rect 13780 14804 13786 14816
rect 13924 14804 13952 14903
rect 15672 14872 15700 14903
rect 15930 14900 15936 14903
rect 15988 14900 15994 14952
rect 17310 14900 17316 14952
rect 17368 14940 17374 14952
rect 17681 14943 17739 14949
rect 17681 14940 17693 14943
rect 17368 14912 17693 14940
rect 17368 14900 17374 14912
rect 17681 14909 17693 14912
rect 17727 14909 17739 14943
rect 17681 14903 17739 14909
rect 17954 14900 17960 14952
rect 18012 14900 18018 14952
rect 18046 14900 18052 14952
rect 18104 14940 18110 14952
rect 18800 14940 18828 14980
rect 19150 14968 19156 14980
rect 19208 14968 19214 15020
rect 19702 14968 19708 15020
rect 19760 14968 19766 15020
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 20349 15011 20407 15017
rect 20349 15008 20361 15011
rect 20027 14980 20361 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 20349 14977 20361 14980
rect 20395 14977 20407 15011
rect 20640 15008 20668 15048
rect 20717 15045 20729 15079
rect 20763 15076 20775 15079
rect 21729 15079 21787 15085
rect 20763 15048 21588 15076
rect 20763 15045 20775 15048
rect 20717 15039 20775 15045
rect 20898 15008 20904 15020
rect 20640 14980 20904 15008
rect 20349 14971 20407 14977
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 21450 14968 21456 15020
rect 21508 14968 21514 15020
rect 18104 14912 18828 14940
rect 19061 14943 19119 14949
rect 18104 14900 18110 14912
rect 19061 14909 19073 14943
rect 19107 14940 19119 14943
rect 19242 14940 19248 14952
rect 19107 14912 19248 14940
rect 19107 14909 19119 14912
rect 19061 14903 19119 14909
rect 19242 14900 19248 14912
rect 19300 14900 19306 14952
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14940 19671 14943
rect 20438 14940 20444 14952
rect 19659 14912 20444 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 20438 14900 20444 14912
rect 20496 14900 20502 14952
rect 20530 14900 20536 14952
rect 20588 14900 20594 14952
rect 21358 14900 21364 14952
rect 21416 14900 21422 14952
rect 21560 14940 21588 15048
rect 21729 15045 21741 15079
rect 21775 15076 21787 15079
rect 22005 15079 22063 15085
rect 22005 15076 22017 15079
rect 21775 15048 22017 15076
rect 21775 15045 21787 15048
rect 21729 15039 21787 15045
rect 22005 15045 22017 15048
rect 22051 15045 22063 15079
rect 22005 15039 22063 15045
rect 21821 15011 21879 15017
rect 21821 14977 21833 15011
rect 21867 15008 21879 15011
rect 22373 15011 22431 15017
rect 22373 15008 22385 15011
rect 21867 14980 22385 15008
rect 21867 14977 21879 14980
rect 21821 14971 21879 14977
rect 22373 14977 22385 14980
rect 22419 14977 22431 15011
rect 22373 14971 22431 14977
rect 21913 14943 21971 14949
rect 21913 14940 21925 14943
rect 21560 14912 21925 14940
rect 21913 14909 21925 14912
rect 21959 14909 21971 14943
rect 21913 14903 21971 14909
rect 22094 14900 22100 14952
rect 22152 14940 22158 14952
rect 22281 14943 22339 14949
rect 22281 14940 22293 14943
rect 22152 14912 22293 14940
rect 22152 14900 22158 14912
rect 22281 14909 22293 14912
rect 22327 14940 22339 14943
rect 22557 14943 22615 14949
rect 22557 14940 22569 14943
rect 22327 14912 22569 14940
rect 22327 14909 22339 14912
rect 22281 14903 22339 14909
rect 22557 14909 22569 14912
rect 22603 14909 22615 14943
rect 22557 14903 22615 14909
rect 22646 14900 22652 14952
rect 22704 14900 22710 14952
rect 16390 14872 16396 14884
rect 15672 14844 16396 14872
rect 15948 14816 15976 14844
rect 16390 14832 16396 14844
rect 16448 14832 16454 14884
rect 17497 14875 17555 14881
rect 17497 14841 17509 14875
rect 17543 14872 17555 14875
rect 17770 14872 17776 14884
rect 17543 14844 17776 14872
rect 17543 14841 17555 14844
rect 17497 14835 17555 14841
rect 17770 14832 17776 14844
rect 17828 14832 17834 14884
rect 18233 14875 18291 14881
rect 18233 14841 18245 14875
rect 18279 14872 18291 14875
rect 18322 14872 18328 14884
rect 18279 14844 18328 14872
rect 18279 14841 18291 14844
rect 18233 14835 18291 14841
rect 18322 14832 18328 14844
rect 18380 14832 18386 14884
rect 19426 14832 19432 14884
rect 19484 14872 19490 14884
rect 20257 14875 20315 14881
rect 20257 14872 20269 14875
rect 19484 14844 20269 14872
rect 19484 14832 19490 14844
rect 20257 14841 20269 14844
rect 20303 14841 20315 14875
rect 20257 14835 20315 14841
rect 22189 14875 22247 14881
rect 22189 14841 22201 14875
rect 22235 14872 22247 14875
rect 22664 14872 22692 14900
rect 22235 14844 22692 14872
rect 22235 14841 22247 14844
rect 22189 14835 22247 14841
rect 13780 14776 13952 14804
rect 13780 14764 13786 14776
rect 15930 14764 15936 14816
rect 15988 14764 15994 14816
rect 22370 14764 22376 14816
rect 22428 14764 22434 14816
rect 552 14714 23368 14736
rect 552 14662 4322 14714
rect 4374 14662 4386 14714
rect 4438 14662 4450 14714
rect 4502 14662 4514 14714
rect 4566 14662 4578 14714
rect 4630 14662 23368 14714
rect 552 14640 23368 14662
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 10008 14572 10149 14600
rect 10008 14560 10014 14572
rect 10137 14569 10149 14572
rect 10183 14600 10195 14603
rect 11057 14603 11115 14609
rect 11057 14600 11069 14603
rect 10183 14572 11069 14600
rect 10183 14569 10195 14572
rect 10137 14563 10195 14569
rect 4246 14492 4252 14544
rect 4304 14532 4310 14544
rect 4494 14535 4552 14541
rect 4494 14532 4506 14535
rect 4304 14504 4506 14532
rect 4304 14492 4310 14504
rect 4494 14501 4506 14504
rect 4540 14501 4552 14535
rect 4494 14495 4552 14501
rect 8018 14492 8024 14544
rect 8076 14532 8082 14544
rect 9585 14535 9643 14541
rect 8076 14504 9352 14532
rect 8076 14492 8082 14504
rect 7190 14464 7196 14476
rect 4264 14436 7196 14464
rect 4264 14405 4292 14436
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 7837 14467 7895 14473
rect 7837 14433 7849 14467
rect 7883 14464 7895 14467
rect 8294 14464 8300 14476
rect 7883 14436 8300 14464
rect 7883 14433 7895 14436
rect 7837 14427 7895 14433
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8390 14467 8448 14473
rect 8390 14433 8402 14467
rect 8436 14433 8448 14467
rect 8390 14427 8448 14433
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 9214 14464 9220 14476
rect 9171 14436 9220 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14396 7987 14399
rect 8110 14396 8116 14408
rect 7975 14368 8116 14396
rect 7975 14365 7987 14368
rect 7929 14359 7987 14365
rect 8110 14356 8116 14368
rect 8168 14396 8174 14408
rect 8404 14396 8432 14427
rect 9214 14424 9220 14436
rect 9272 14424 9278 14476
rect 9324 14473 9352 14504
rect 9585 14501 9597 14535
rect 9631 14532 9643 14535
rect 9674 14532 9680 14544
rect 9631 14504 9680 14532
rect 9631 14501 9643 14504
rect 9585 14495 9643 14501
rect 9674 14492 9680 14504
rect 9732 14532 9738 14544
rect 10226 14532 10232 14544
rect 9732 14504 10232 14532
rect 9732 14492 9738 14504
rect 10226 14492 10232 14504
rect 10284 14492 10290 14544
rect 10318 14492 10324 14544
rect 10376 14532 10382 14544
rect 10594 14541 10600 14544
rect 10565 14535 10600 14541
rect 10565 14532 10577 14535
rect 10376 14504 10577 14532
rect 10376 14492 10382 14504
rect 10565 14501 10577 14504
rect 10565 14495 10600 14501
rect 10594 14492 10600 14495
rect 10652 14492 10658 14544
rect 10796 14541 10824 14572
rect 11057 14569 11069 14572
rect 11103 14569 11115 14603
rect 11057 14563 11115 14569
rect 11422 14560 11428 14612
rect 11480 14600 11486 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 11480 14572 13001 14600
rect 11480 14560 11486 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 13633 14603 13691 14609
rect 13633 14569 13645 14603
rect 13679 14600 13691 14603
rect 14458 14600 14464 14612
rect 13679 14572 14464 14600
rect 13679 14569 13691 14572
rect 13633 14563 13691 14569
rect 14458 14560 14464 14572
rect 14516 14560 14522 14612
rect 17310 14560 17316 14612
rect 17368 14600 17374 14612
rect 17497 14603 17555 14609
rect 17497 14600 17509 14603
rect 17368 14572 17509 14600
rect 17368 14560 17374 14572
rect 17497 14569 17509 14572
rect 17543 14569 17555 14603
rect 17497 14563 17555 14569
rect 17681 14603 17739 14609
rect 17681 14569 17693 14603
rect 17727 14600 17739 14603
rect 17954 14600 17960 14612
rect 17727 14572 17960 14600
rect 17727 14569 17739 14572
rect 17681 14563 17739 14569
rect 10755 14535 10824 14541
rect 10755 14501 10767 14535
rect 10801 14504 10824 14535
rect 13817 14535 13875 14541
rect 13817 14532 13829 14535
rect 12912 14504 13829 14532
rect 10801 14501 10813 14504
rect 10755 14495 10813 14501
rect 9309 14467 9367 14473
rect 9309 14433 9321 14467
rect 9355 14433 9367 14467
rect 9309 14427 9367 14433
rect 9769 14467 9827 14473
rect 9769 14433 9781 14467
rect 9815 14464 9827 14467
rect 9858 14464 9864 14476
rect 9815 14436 9864 14464
rect 9815 14433 9827 14436
rect 9769 14427 9827 14433
rect 8168 14368 8432 14396
rect 8168 14356 8174 14368
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 9784 14396 9812 14427
rect 9858 14424 9864 14436
rect 9916 14424 9922 14476
rect 10042 14424 10048 14476
rect 10100 14464 10106 14476
rect 10965 14467 11023 14473
rect 10965 14464 10977 14467
rect 10100 14436 10977 14464
rect 10100 14424 10106 14436
rect 9640 14368 9812 14396
rect 9640 14356 9646 14368
rect 8665 14331 8723 14337
rect 8665 14297 8677 14331
rect 8711 14328 8723 14331
rect 8938 14328 8944 14340
rect 8711 14300 8944 14328
rect 8711 14297 8723 14300
rect 8665 14291 8723 14297
rect 8938 14288 8944 14300
rect 8996 14288 9002 14340
rect 9858 14288 9864 14340
rect 9916 14328 9922 14340
rect 10321 14331 10379 14337
rect 10321 14328 10333 14331
rect 9916 14300 10333 14328
rect 9916 14288 9922 14300
rect 10321 14297 10333 14300
rect 10367 14297 10379 14331
rect 10321 14291 10379 14297
rect 5626 14220 5632 14272
rect 5684 14220 5690 14272
rect 8205 14263 8263 14269
rect 8205 14229 8217 14263
rect 8251 14260 8263 14263
rect 8386 14260 8392 14272
rect 8251 14232 8392 14260
rect 8251 14229 8263 14232
rect 8205 14223 8263 14229
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 9217 14263 9275 14269
rect 9217 14229 9229 14263
rect 9263 14260 9275 14263
rect 9766 14260 9772 14272
rect 9263 14232 9772 14260
rect 9263 14229 9275 14232
rect 9217 14223 9275 14229
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 9950 14220 9956 14272
rect 10008 14220 10014 14272
rect 10134 14220 10140 14272
rect 10192 14260 10198 14272
rect 10410 14260 10416 14272
rect 10192 14232 10416 14260
rect 10192 14220 10198 14232
rect 10410 14220 10416 14232
rect 10468 14220 10474 14272
rect 10580 14269 10608 14436
rect 10965 14433 10977 14436
rect 11011 14433 11023 14467
rect 10965 14427 11023 14433
rect 11241 14467 11299 14473
rect 11241 14433 11253 14467
rect 11287 14433 11299 14467
rect 11241 14427 11299 14433
rect 10686 14356 10692 14408
rect 10744 14396 10750 14408
rect 11256 14396 11284 14427
rect 12066 14424 12072 14476
rect 12124 14464 12130 14476
rect 12912 14473 12940 14504
rect 13817 14501 13829 14504
rect 13863 14501 13875 14535
rect 13817 14495 13875 14501
rect 16384 14535 16442 14541
rect 16384 14501 16396 14535
rect 16430 14532 16442 14535
rect 16758 14532 16764 14544
rect 16430 14504 16764 14532
rect 16430 14501 16442 14504
rect 16384 14495 16442 14501
rect 16758 14492 16764 14504
rect 16816 14492 16822 14544
rect 12897 14467 12955 14473
rect 12897 14464 12909 14467
rect 12124 14436 12909 14464
rect 12124 14424 12130 14436
rect 12897 14433 12909 14436
rect 12943 14433 12955 14467
rect 12897 14427 12955 14433
rect 13170 14424 13176 14476
rect 13228 14424 13234 14476
rect 13357 14467 13415 14473
rect 13357 14433 13369 14467
rect 13403 14464 13415 14467
rect 13538 14464 13544 14476
rect 13403 14436 13544 14464
rect 13403 14433 13415 14436
rect 13357 14427 13415 14433
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 13722 14424 13728 14476
rect 13780 14424 13786 14476
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 14001 14467 14059 14473
rect 14001 14464 14013 14467
rect 13964 14436 14013 14464
rect 13964 14424 13970 14436
rect 14001 14433 14013 14436
rect 14047 14433 14059 14467
rect 17512 14464 17540 14563
rect 17954 14560 17960 14572
rect 18012 14600 18018 14612
rect 18065 14603 18123 14609
rect 18065 14600 18077 14603
rect 18012 14572 18077 14600
rect 18012 14560 18018 14572
rect 18065 14569 18077 14572
rect 18111 14569 18123 14603
rect 18065 14563 18123 14569
rect 19426 14560 19432 14612
rect 19484 14560 19490 14612
rect 21818 14600 21824 14612
rect 21284 14572 21824 14600
rect 17865 14535 17923 14541
rect 17865 14501 17877 14535
rect 17911 14532 17923 14535
rect 18322 14532 18328 14544
rect 17911 14504 18328 14532
rect 17911 14501 17923 14504
rect 17865 14495 17923 14501
rect 18322 14492 18328 14504
rect 18380 14492 18386 14544
rect 17589 14467 17647 14473
rect 17589 14464 17601 14467
rect 17512 14436 17601 14464
rect 14001 14427 14059 14433
rect 17589 14433 17601 14436
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 17770 14424 17776 14476
rect 17828 14424 17834 14476
rect 18506 14424 18512 14476
rect 18564 14424 18570 14476
rect 18966 14424 18972 14476
rect 19024 14424 19030 14476
rect 21284 14473 21312 14572
rect 21818 14560 21824 14572
rect 21876 14560 21882 14612
rect 22830 14560 22836 14612
rect 22888 14600 22894 14612
rect 23017 14603 23075 14609
rect 23017 14600 23029 14603
rect 22888 14572 23029 14600
rect 22888 14560 22894 14572
rect 23017 14569 23029 14572
rect 23063 14569 23075 14603
rect 23017 14563 23075 14569
rect 21637 14535 21695 14541
rect 21637 14501 21649 14535
rect 21683 14532 21695 14535
rect 21683 14504 22876 14532
rect 21683 14501 21695 14504
rect 21637 14495 21695 14501
rect 19245 14467 19303 14473
rect 19245 14433 19257 14467
rect 19291 14433 19303 14467
rect 19245 14427 19303 14433
rect 21269 14467 21327 14473
rect 21269 14433 21281 14467
rect 21315 14433 21327 14467
rect 21269 14427 21327 14433
rect 21361 14467 21419 14473
rect 21361 14433 21373 14467
rect 21407 14433 21419 14467
rect 21361 14427 21419 14433
rect 21545 14467 21603 14473
rect 21545 14433 21557 14467
rect 21591 14464 21603 14467
rect 21726 14464 21732 14476
rect 21591 14436 21732 14464
rect 21591 14433 21603 14436
rect 21545 14427 21603 14433
rect 10744 14368 11284 14396
rect 10744 14356 10750 14368
rect 13262 14356 13268 14408
rect 13320 14396 13326 14408
rect 13924 14396 13952 14424
rect 13320 14368 13952 14396
rect 13320 14356 13326 14368
rect 15930 14356 15936 14408
rect 15988 14396 15994 14408
rect 16117 14399 16175 14405
rect 16117 14396 16129 14399
rect 15988 14368 16129 14396
rect 15988 14356 15994 14368
rect 16117 14365 16129 14368
rect 16163 14365 16175 14399
rect 16117 14359 16175 14365
rect 18598 14356 18604 14408
rect 18656 14356 18662 14408
rect 18782 14356 18788 14408
rect 18840 14396 18846 14408
rect 19061 14399 19119 14405
rect 19061 14396 19073 14399
rect 18840 14368 19073 14396
rect 18840 14356 18846 14368
rect 19061 14365 19073 14368
rect 19107 14365 19119 14399
rect 19061 14359 19119 14365
rect 18877 14331 18935 14337
rect 18877 14297 18889 14331
rect 18923 14328 18935 14331
rect 19260 14328 19288 14427
rect 21376 14396 21404 14427
rect 21726 14424 21732 14436
rect 21784 14424 21790 14476
rect 21818 14424 21824 14476
rect 21876 14424 21882 14476
rect 21913 14467 21971 14473
rect 21913 14433 21925 14467
rect 21959 14433 21971 14467
rect 21913 14427 21971 14433
rect 21634 14396 21640 14408
rect 21376 14368 21640 14396
rect 21634 14356 21640 14368
rect 21692 14396 21698 14408
rect 21928 14396 21956 14427
rect 22002 14424 22008 14476
rect 22060 14424 22066 14476
rect 22186 14473 22192 14476
rect 22143 14467 22192 14473
rect 22143 14433 22155 14467
rect 22189 14433 22192 14467
rect 22143 14427 22192 14433
rect 22186 14424 22192 14427
rect 22244 14424 22250 14476
rect 22373 14467 22431 14473
rect 22373 14433 22385 14467
rect 22419 14464 22431 14467
rect 22462 14464 22468 14476
rect 22419 14436 22468 14464
rect 22419 14433 22431 14436
rect 22373 14427 22431 14433
rect 22462 14424 22468 14436
rect 22520 14424 22526 14476
rect 22848 14473 22876 14504
rect 22833 14467 22891 14473
rect 22833 14433 22845 14467
rect 22879 14433 22891 14467
rect 22833 14427 22891 14433
rect 21692 14368 21956 14396
rect 21692 14356 21698 14368
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 22554 14396 22560 14408
rect 22336 14368 22560 14396
rect 22336 14356 22342 14368
rect 22554 14356 22560 14368
rect 22612 14356 22618 14408
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14365 22707 14399
rect 22649 14359 22707 14365
rect 18923 14300 19288 14328
rect 21545 14331 21603 14337
rect 18923 14297 18935 14300
rect 18877 14291 18935 14297
rect 21545 14297 21557 14331
rect 21591 14328 21603 14331
rect 22664 14328 22692 14359
rect 21591 14300 22692 14328
rect 21591 14297 21603 14300
rect 21545 14291 21603 14297
rect 10575 14263 10633 14269
rect 10575 14229 10587 14263
rect 10621 14229 10633 14263
rect 10575 14223 10633 14229
rect 11425 14263 11483 14269
rect 11425 14229 11437 14263
rect 11471 14260 11483 14263
rect 12710 14260 12716 14272
rect 11471 14232 12716 14260
rect 11471 14229 11483 14232
rect 11425 14223 11483 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14185 14263 14243 14269
rect 14185 14260 14197 14263
rect 13872 14232 14197 14260
rect 13872 14220 13878 14232
rect 14185 14229 14197 14232
rect 14231 14229 14243 14263
rect 14185 14223 14243 14229
rect 18046 14220 18052 14272
rect 18104 14220 18110 14272
rect 18230 14220 18236 14272
rect 18288 14220 18294 14272
rect 19058 14220 19064 14272
rect 19116 14220 19122 14272
rect 22370 14220 22376 14272
rect 22428 14260 22434 14272
rect 22465 14263 22523 14269
rect 22465 14260 22477 14263
rect 22428 14232 22477 14260
rect 22428 14220 22434 14232
rect 22465 14229 22477 14232
rect 22511 14229 22523 14263
rect 22465 14223 22523 14229
rect 552 14170 23368 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 23368 14170
rect 552 14096 23368 14118
rect 4157 14059 4215 14065
rect 4157 14025 4169 14059
rect 4203 14056 4215 14059
rect 5166 14056 5172 14068
rect 4203 14028 5172 14056
rect 4203 14025 4215 14028
rect 4157 14019 4215 14025
rect 5166 14016 5172 14028
rect 5224 14056 5230 14068
rect 5224 14028 6132 14056
rect 5224 14016 5230 14028
rect 5629 13991 5687 13997
rect 5629 13957 5641 13991
rect 5675 13957 5687 13991
rect 5629 13951 5687 13957
rect 5644 13920 5672 13951
rect 6104 13929 6132 14028
rect 9030 14016 9036 14068
rect 9088 14056 9094 14068
rect 9582 14056 9588 14068
rect 9088 14028 9588 14056
rect 9088 14016 9094 14028
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 10410 14056 10416 14068
rect 9876 14028 10416 14056
rect 8573 13991 8631 13997
rect 8573 13957 8585 13991
rect 8619 13988 8631 13991
rect 9214 13988 9220 14000
rect 8619 13960 9220 13988
rect 8619 13957 8631 13960
rect 8573 13951 8631 13957
rect 9214 13948 9220 13960
rect 9272 13948 9278 14000
rect 9876 13997 9904 14028
rect 10410 14016 10416 14028
rect 10468 14056 10474 14068
rect 10873 14059 10931 14065
rect 10873 14056 10885 14059
rect 10468 14028 10885 14056
rect 10468 14016 10474 14028
rect 10873 14025 10885 14028
rect 10919 14025 10931 14059
rect 10873 14019 10931 14025
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 12492 14028 12664 14056
rect 12492 14016 12498 14028
rect 9861 13991 9919 13997
rect 9861 13957 9873 13991
rect 9907 13957 9919 13991
rect 9861 13951 9919 13957
rect 11057 13991 11115 13997
rect 11057 13957 11069 13991
rect 11103 13957 11115 13991
rect 11057 13951 11115 13957
rect 12161 13991 12219 13997
rect 12161 13957 12173 13991
rect 12207 13988 12219 13991
rect 12526 13988 12532 14000
rect 12207 13960 12532 13988
rect 12207 13957 12219 13960
rect 12161 13951 12219 13957
rect 5460 13892 5672 13920
rect 6089 13923 6147 13929
rect 5281 13855 5339 13861
rect 5281 13821 5293 13855
rect 5327 13852 5339 13855
rect 5460 13852 5488 13892
rect 6089 13889 6101 13923
rect 6135 13889 6147 13923
rect 6089 13883 6147 13889
rect 6273 13923 6331 13929
rect 6273 13889 6285 13923
rect 6319 13920 6331 13923
rect 6914 13920 6920 13932
rect 6319 13892 6920 13920
rect 6319 13889 6331 13892
rect 6273 13883 6331 13889
rect 6914 13880 6920 13892
rect 6972 13920 6978 13932
rect 8110 13920 8116 13932
rect 6972 13892 8116 13920
rect 6972 13880 6978 13892
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 8996 13892 9720 13920
rect 8996 13880 9002 13892
rect 5327 13824 5488 13852
rect 5537 13855 5595 13861
rect 5327 13821 5339 13824
rect 5281 13815 5339 13821
rect 5537 13821 5549 13855
rect 5583 13852 5595 13855
rect 7190 13852 7196 13864
rect 5583 13824 7196 13852
rect 5583 13821 5595 13824
rect 5537 13815 5595 13821
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 8386 13812 8392 13864
rect 8444 13812 8450 13864
rect 8570 13812 8576 13864
rect 8628 13852 8634 13864
rect 8754 13852 8760 13864
rect 8628 13824 8760 13852
rect 8628 13812 8634 13824
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 9030 13852 9036 13864
rect 8956 13824 9036 13852
rect 5442 13744 5448 13796
rect 5500 13784 5506 13796
rect 8956 13793 8984 13824
rect 9030 13812 9036 13824
rect 9088 13812 9094 13864
rect 9692 13861 9720 13892
rect 9766 13880 9772 13932
rect 9824 13920 9830 13932
rect 11072 13920 11100 13951
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 11149 13923 11207 13929
rect 11149 13920 11161 13923
rect 9824 13892 10456 13920
rect 11072 13892 11161 13920
rect 9824 13880 9830 13892
rect 9125 13855 9183 13861
rect 9125 13821 9137 13855
rect 9171 13852 9183 13855
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 9171 13824 9505 13852
rect 9171 13821 9183 13824
rect 9125 13815 9183 13821
rect 9493 13821 9505 13824
rect 9539 13852 9551 13855
rect 9677 13855 9735 13861
rect 9539 13824 9628 13852
rect 9539 13821 9551 13824
rect 9493 13815 9551 13821
rect 9600 13796 9628 13824
rect 9677 13821 9689 13855
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 9858 13812 9864 13864
rect 9916 13852 9922 13864
rect 9953 13855 10011 13861
rect 9953 13852 9965 13855
rect 9916 13824 9965 13852
rect 9916 13812 9922 13824
rect 9953 13821 9965 13824
rect 9999 13821 10011 13855
rect 9953 13815 10011 13821
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13852 10103 13855
rect 10134 13852 10140 13864
rect 10091 13824 10140 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 10318 13812 10324 13864
rect 10376 13812 10382 13864
rect 10428 13861 10456 13892
rect 11149 13889 11161 13892
rect 11195 13889 11207 13923
rect 11149 13883 11207 13889
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13920 12403 13923
rect 12434 13920 12440 13932
rect 12391 13892 12440 13920
rect 12391 13889 12403 13892
rect 12345 13883 12403 13889
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 12636 13929 12664 14028
rect 13814 14016 13820 14068
rect 13872 14016 13878 14068
rect 14185 14059 14243 14065
rect 14185 14056 14197 14059
rect 13924 14028 14197 14056
rect 13357 13991 13415 13997
rect 13357 13957 13369 13991
rect 13403 13988 13415 13991
rect 13924 13988 13952 14028
rect 14185 14025 14197 14028
rect 14231 14025 14243 14059
rect 14185 14019 14243 14025
rect 16758 14016 16764 14068
rect 16816 14056 16822 14068
rect 17405 14059 17463 14065
rect 17405 14056 17417 14059
rect 16816 14028 17417 14056
rect 16816 14016 16822 14028
rect 17405 14025 17417 14028
rect 17451 14025 17463 14059
rect 17405 14019 17463 14025
rect 17589 14059 17647 14065
rect 17589 14025 17601 14059
rect 17635 14056 17647 14059
rect 18046 14056 18052 14068
rect 17635 14028 18052 14056
rect 17635 14025 17647 14028
rect 17589 14019 17647 14025
rect 13403 13960 13952 13988
rect 14001 13991 14059 13997
rect 13403 13957 13415 13960
rect 13357 13951 13415 13957
rect 14001 13957 14013 13991
rect 14047 13957 14059 13991
rect 14001 13951 14059 13957
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13889 12679 13923
rect 12621 13883 12679 13889
rect 12710 13880 12716 13932
rect 12768 13880 12774 13932
rect 12802 13880 12808 13932
rect 12860 13880 12866 13932
rect 13814 13920 13820 13932
rect 13096 13892 13820 13920
rect 10413 13855 10471 13861
rect 10413 13821 10425 13855
rect 10459 13852 10471 13855
rect 10459 13827 10932 13852
rect 10459 13824 10977 13827
rect 10459 13821 10471 13824
rect 10413 13815 10471 13821
rect 10904 13821 10977 13824
rect 5997 13787 6055 13793
rect 5997 13784 6009 13787
rect 5500 13756 6009 13784
rect 5500 13744 5506 13756
rect 5997 13753 6009 13756
rect 6043 13753 6055 13787
rect 5997 13747 6055 13753
rect 8941 13787 8999 13793
rect 8941 13753 8953 13787
rect 8987 13753 8999 13787
rect 8941 13747 8999 13753
rect 9217 13787 9275 13793
rect 9217 13753 9229 13787
rect 9263 13753 9275 13787
rect 9217 13747 9275 13753
rect 8754 13676 8760 13728
rect 8812 13676 8818 13728
rect 9232 13716 9260 13747
rect 9582 13744 9588 13796
rect 9640 13744 9646 13796
rect 10229 13787 10287 13793
rect 10229 13753 10241 13787
rect 10275 13753 10287 13787
rect 10689 13787 10747 13793
rect 10904 13790 10931 13821
rect 10689 13784 10701 13787
rect 10229 13747 10287 13753
rect 10428 13756 10701 13784
rect 10134 13716 10140 13728
rect 9232 13688 10140 13716
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 10244 13716 10272 13747
rect 10428 13728 10456 13756
rect 10689 13753 10701 13756
rect 10735 13753 10747 13787
rect 10919 13787 10931 13790
rect 10965 13787 10977 13821
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11333 13855 11391 13861
rect 11333 13852 11345 13855
rect 11112 13824 11345 13852
rect 11112 13812 11118 13824
rect 11333 13821 11345 13824
rect 11379 13821 11391 13855
rect 11333 13815 11391 13821
rect 11422 13812 11428 13864
rect 11480 13812 11486 13864
rect 12066 13812 12072 13864
rect 12124 13812 12130 13864
rect 13096 13861 13124 13892
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 12253 13855 12311 13861
rect 12253 13821 12265 13855
rect 12299 13852 12311 13855
rect 12529 13855 12587 13861
rect 12299 13824 12434 13852
rect 12299 13821 12311 13824
rect 12253 13815 12311 13821
rect 10919 13781 10977 13787
rect 10689 13747 10747 13753
rect 10410 13716 10416 13728
rect 10244 13688 10416 13716
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 10597 13719 10655 13725
rect 10597 13685 10609 13719
rect 10643 13716 10655 13719
rect 11054 13716 11060 13728
rect 10643 13688 11060 13716
rect 10643 13685 10655 13688
rect 10597 13679 10655 13685
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 11146 13676 11152 13728
rect 11204 13676 11210 13728
rect 12406 13716 12434 13824
rect 12529 13821 12541 13855
rect 12575 13821 12587 13855
rect 12529 13815 12587 13821
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 12544 13784 12572 13815
rect 13170 13812 13176 13864
rect 13228 13812 13234 13864
rect 13357 13855 13415 13861
rect 13357 13821 13369 13855
rect 13403 13852 13415 13855
rect 13538 13852 13544 13864
rect 13403 13824 13544 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 13538 13812 13544 13824
rect 13596 13852 13602 13864
rect 14016 13852 14044 13951
rect 14090 13948 14096 14000
rect 14148 13988 14154 14000
rect 14277 13991 14335 13997
rect 14277 13988 14289 13991
rect 14148 13960 14289 13988
rect 14148 13948 14154 13960
rect 14277 13957 14289 13960
rect 14323 13957 14335 13991
rect 17420 13988 17448 14019
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 19058 14016 19064 14068
rect 19116 14016 19122 14068
rect 21266 14056 21272 14068
rect 20364 14028 21272 14056
rect 17770 13988 17776 14000
rect 17420 13960 17776 13988
rect 14277 13951 14335 13957
rect 17770 13948 17776 13960
rect 17828 13948 17834 14000
rect 17954 13948 17960 14000
rect 18012 13948 18018 14000
rect 14366 13880 14372 13932
rect 14424 13920 14430 13932
rect 15381 13923 15439 13929
rect 15381 13920 15393 13923
rect 14424 13892 15393 13920
rect 14424 13880 14430 13892
rect 15381 13889 15393 13892
rect 15427 13920 15439 13923
rect 17126 13920 17132 13932
rect 15427 13892 17132 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 20364 13929 20392 14028
rect 21266 14016 21272 14028
rect 21324 14056 21330 14068
rect 21542 14056 21548 14068
rect 21324 14028 21548 14056
rect 21324 14016 21330 14028
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 22830 13988 22836 14000
rect 22066 13960 22836 13988
rect 20349 13923 20407 13929
rect 17236 13892 18000 13920
rect 14093 13855 14151 13861
rect 14093 13852 14105 13855
rect 13596 13827 13876 13852
rect 13596 13824 13921 13827
rect 14016 13824 14105 13852
rect 13596 13812 13602 13824
rect 13848 13821 13921 13824
rect 12618 13784 12624 13796
rect 12544 13756 12624 13784
rect 12618 13744 12624 13756
rect 12676 13784 12682 13796
rect 13188 13784 13216 13812
rect 12676 13756 13216 13784
rect 12676 13744 12682 13756
rect 13630 13744 13636 13796
rect 13688 13744 13694 13796
rect 13848 13790 13875 13821
rect 13863 13787 13875 13790
rect 13909 13787 13921 13821
rect 14093 13821 14105 13824
rect 14139 13821 14151 13855
rect 14093 13815 14151 13821
rect 15286 13812 15292 13864
rect 15344 13852 15350 13864
rect 15565 13855 15623 13861
rect 15565 13852 15577 13855
rect 15344 13824 15577 13852
rect 15344 13812 15350 13824
rect 15565 13821 15577 13824
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 17236 13796 17264 13892
rect 17681 13855 17739 13861
rect 17681 13821 17693 13855
rect 17727 13821 17739 13855
rect 17681 13815 17739 13821
rect 13863 13781 13921 13787
rect 15470 13744 15476 13796
rect 15528 13784 15534 13796
rect 15657 13787 15715 13793
rect 15657 13784 15669 13787
rect 15528 13756 15669 13784
rect 15528 13744 15534 13756
rect 15657 13753 15669 13756
rect 15703 13753 15715 13787
rect 15657 13747 15715 13753
rect 17218 13744 17224 13796
rect 17276 13744 17282 13796
rect 12802 13716 12808 13728
rect 12406 13688 12808 13716
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 13173 13719 13231 13725
rect 13173 13685 13185 13719
rect 13219 13716 13231 13719
rect 13648 13716 13676 13744
rect 13219 13688 13676 13716
rect 13219 13685 13231 13688
rect 13173 13679 13231 13685
rect 16022 13676 16028 13728
rect 16080 13676 16086 13728
rect 17126 13676 17132 13728
rect 17184 13716 17190 13728
rect 17421 13719 17479 13725
rect 17421 13716 17433 13719
rect 17184 13688 17433 13716
rect 17184 13676 17190 13688
rect 17421 13685 17433 13688
rect 17467 13716 17479 13719
rect 17696 13716 17724 13815
rect 17770 13812 17776 13864
rect 17828 13812 17834 13864
rect 17972 13861 18000 13892
rect 20349 13889 20361 13923
rect 20395 13889 20407 13923
rect 22066 13920 22094 13960
rect 22830 13948 22836 13960
rect 22888 13948 22894 14000
rect 20349 13883 20407 13889
rect 22020 13892 22094 13920
rect 22189 13923 22247 13929
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13821 18015 13855
rect 17957 13815 18015 13821
rect 18230 13812 18236 13864
rect 18288 13852 18294 13864
rect 18877 13855 18935 13861
rect 18877 13852 18889 13855
rect 18288 13824 18889 13852
rect 18288 13812 18294 13824
rect 18877 13821 18889 13824
rect 18923 13821 18935 13855
rect 18877 13815 18935 13821
rect 20616 13855 20674 13861
rect 20616 13821 20628 13855
rect 20662 13852 20674 13855
rect 20898 13852 20904 13864
rect 20662 13824 20904 13852
rect 20662 13821 20674 13824
rect 20616 13815 20674 13821
rect 20898 13812 20904 13824
rect 20956 13812 20962 13864
rect 22020 13861 22048 13892
rect 22189 13889 22201 13923
rect 22235 13920 22247 13923
rect 22738 13920 22744 13932
rect 22235 13892 22744 13920
rect 22235 13889 22247 13892
rect 22189 13883 22247 13889
rect 22738 13880 22744 13892
rect 22796 13880 22802 13932
rect 22005 13855 22063 13861
rect 22005 13821 22017 13855
rect 22051 13821 22063 13855
rect 22005 13815 22063 13821
rect 18690 13744 18696 13796
rect 18748 13744 18754 13796
rect 17467 13688 17724 13716
rect 17467 13685 17479 13688
rect 17421 13679 17479 13685
rect 21358 13676 21364 13728
rect 21416 13716 21422 13728
rect 21729 13719 21787 13725
rect 21729 13716 21741 13719
rect 21416 13688 21741 13716
rect 21416 13676 21422 13688
rect 21729 13685 21741 13688
rect 21775 13685 21787 13719
rect 21729 13679 21787 13685
rect 21818 13676 21824 13728
rect 21876 13676 21882 13728
rect 552 13626 23368 13648
rect 552 13574 4322 13626
rect 4374 13574 4386 13626
rect 4438 13574 4450 13626
rect 4502 13574 4514 13626
rect 4566 13574 4578 13626
rect 4630 13574 23368 13626
rect 552 13552 23368 13574
rect 5350 13472 5356 13524
rect 5408 13472 5414 13524
rect 6273 13515 6331 13521
rect 6273 13481 6285 13515
rect 6319 13512 6331 13515
rect 6362 13512 6368 13524
rect 6319 13484 6368 13512
rect 6319 13481 6331 13484
rect 6273 13475 6331 13481
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 8297 13515 8355 13521
rect 8297 13481 8309 13515
rect 8343 13512 8355 13515
rect 8386 13512 8392 13524
rect 8343 13484 8392 13512
rect 8343 13481 8355 13484
rect 8297 13475 8355 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 10410 13472 10416 13524
rect 10468 13472 10474 13524
rect 12437 13515 12495 13521
rect 12437 13481 12449 13515
rect 12483 13512 12495 13515
rect 12710 13512 12716 13524
rect 12483 13484 12716 13512
rect 12483 13481 12495 13484
rect 12437 13475 12495 13481
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 13722 13512 13728 13524
rect 12860 13484 13728 13512
rect 12860 13472 12866 13484
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 14553 13515 14611 13521
rect 14553 13481 14565 13515
rect 14599 13512 14611 13515
rect 15470 13512 15476 13524
rect 14599 13484 15476 13512
rect 14599 13481 14611 13484
rect 14553 13475 14611 13481
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 16758 13472 16764 13524
rect 16816 13472 16822 13524
rect 17126 13472 17132 13524
rect 17184 13472 17190 13524
rect 18141 13515 18199 13521
rect 18141 13481 18153 13515
rect 18187 13512 18199 13515
rect 18782 13512 18788 13524
rect 18187 13484 18788 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 18782 13472 18788 13484
rect 18840 13472 18846 13524
rect 21726 13472 21732 13524
rect 21784 13512 21790 13524
rect 22373 13515 22431 13521
rect 22373 13512 22385 13515
rect 21784 13484 22385 13512
rect 21784 13472 21790 13484
rect 22373 13481 22385 13484
rect 22419 13512 22431 13515
rect 22419 13484 22508 13512
rect 22419 13481 22431 13484
rect 22373 13475 22431 13481
rect 8110 13404 8116 13456
rect 8168 13444 8174 13456
rect 8478 13444 8484 13456
rect 8168 13416 8484 13444
rect 8168 13404 8174 13416
rect 8478 13404 8484 13416
rect 8536 13404 8542 13456
rect 8754 13404 8760 13456
rect 8812 13444 8818 13456
rect 10428 13444 10456 13472
rect 8812 13416 9260 13444
rect 8812 13404 8818 13416
rect 5258 13336 5264 13388
rect 5316 13336 5322 13388
rect 6178 13336 6184 13388
rect 6236 13336 6242 13388
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 8570 13376 8576 13388
rect 8435 13348 8576 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 8570 13336 8576 13348
rect 8628 13336 8634 13388
rect 8938 13336 8944 13388
rect 8996 13336 9002 13388
rect 9232 13385 9260 13416
rect 10152 13416 10456 13444
rect 9217 13379 9275 13385
rect 9217 13345 9229 13379
rect 9263 13345 9275 13379
rect 9217 13339 9275 13345
rect 9401 13379 9459 13385
rect 9401 13345 9413 13379
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 5537 13311 5595 13317
rect 5537 13277 5549 13311
rect 5583 13308 5595 13311
rect 6365 13311 6423 13317
rect 6365 13308 6377 13311
rect 5583 13280 6377 13308
rect 5583 13277 5595 13280
rect 5537 13271 5595 13277
rect 6365 13277 6377 13280
rect 6411 13308 6423 13311
rect 6822 13308 6828 13320
rect 6411 13280 6828 13308
rect 6411 13277 6423 13280
rect 6365 13271 6423 13277
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 8956 13308 8984 13336
rect 9416 13308 9444 13339
rect 9950 13336 9956 13388
rect 10008 13336 10014 13388
rect 10152 13385 10180 13416
rect 12526 13404 12532 13456
rect 12584 13444 12590 13456
rect 12584 13416 13124 13444
rect 12584 13404 12590 13416
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 10226 13336 10232 13388
rect 10284 13336 10290 13388
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13345 10471 13379
rect 10413 13339 10471 13345
rect 8956 13280 9444 13308
rect 10042 13268 10048 13320
rect 10100 13308 10106 13320
rect 10428 13308 10456 13339
rect 12342 13336 12348 13388
rect 12400 13336 12406 13388
rect 12618 13336 12624 13388
rect 12676 13336 12682 13388
rect 13096 13385 13124 13416
rect 13262 13385 13268 13388
rect 13081 13379 13139 13385
rect 13081 13345 13093 13379
rect 13127 13345 13139 13379
rect 13081 13339 13139 13345
rect 13235 13379 13268 13385
rect 13235 13345 13247 13379
rect 13235 13339 13268 13345
rect 13262 13336 13268 13339
rect 13320 13336 13326 13388
rect 13814 13336 13820 13388
rect 13872 13336 13878 13388
rect 13909 13379 13967 13385
rect 13909 13345 13921 13379
rect 13955 13376 13967 13379
rect 14366 13376 14372 13388
rect 13955 13348 14372 13376
rect 13955 13345 13967 13348
rect 13909 13339 13967 13345
rect 14366 13336 14372 13348
rect 14424 13336 14430 13388
rect 15488 13376 15516 13472
rect 15688 13447 15746 13453
rect 15688 13413 15700 13447
rect 15734 13444 15746 13447
rect 16022 13444 16028 13456
rect 15734 13416 16028 13444
rect 15734 13413 15746 13416
rect 15688 13407 15746 13413
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 17957 13447 18015 13453
rect 16316 13416 16896 13444
rect 15488 13348 16068 13376
rect 10100 13280 10456 13308
rect 13449 13311 13507 13317
rect 10100 13268 10106 13280
rect 13449 13277 13461 13311
rect 13495 13308 13507 13311
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 13495 13280 13737 13308
rect 13495 13277 13507 13280
rect 13449 13271 13507 13277
rect 13725 13277 13737 13280
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 13998 13268 14004 13320
rect 14056 13268 14062 13320
rect 15930 13268 15936 13320
rect 15988 13268 15994 13320
rect 16040 13308 16068 13348
rect 16316 13320 16344 13416
rect 16390 13336 16396 13388
rect 16448 13376 16454 13388
rect 16868 13385 16896 13416
rect 17957 13413 17969 13447
rect 18003 13444 18015 13447
rect 18046 13444 18052 13456
rect 18003 13416 18052 13444
rect 18003 13413 18015 13416
rect 17957 13407 18015 13413
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 18233 13447 18291 13453
rect 18233 13413 18245 13447
rect 18279 13413 18291 13447
rect 18233 13407 18291 13413
rect 16853 13379 16911 13385
rect 16448 13348 16620 13376
rect 16448 13336 16454 13348
rect 16298 13308 16304 13320
rect 16040 13280 16304 13308
rect 16298 13268 16304 13280
rect 16356 13308 16362 13320
rect 16485 13311 16543 13317
rect 16485 13308 16497 13311
rect 16356 13280 16497 13308
rect 16356 13268 16362 13280
rect 16485 13277 16497 13280
rect 16531 13277 16543 13311
rect 16592 13308 16620 13348
rect 16853 13345 16865 13379
rect 16899 13345 16911 13379
rect 16853 13339 16911 13345
rect 17773 13379 17831 13385
rect 17773 13345 17785 13379
rect 17819 13376 17831 13379
rect 17862 13376 17868 13388
rect 17819 13348 17868 13376
rect 17819 13345 17831 13348
rect 17773 13339 17831 13345
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18248 13376 18276 13407
rect 18414 13404 18420 13456
rect 18472 13453 18478 13456
rect 18472 13447 18491 13453
rect 18479 13413 18491 13447
rect 18472 13407 18491 13413
rect 19797 13447 19855 13453
rect 19797 13413 19809 13447
rect 19843 13444 19855 13447
rect 20806 13444 20812 13456
rect 19843 13416 20812 13444
rect 19843 13413 19855 13416
rect 19797 13407 19855 13413
rect 18472 13404 18478 13407
rect 18322 13376 18328 13388
rect 18248 13348 18328 13376
rect 18322 13336 18328 13348
rect 18380 13376 18386 13388
rect 19150 13376 19156 13388
rect 18380 13348 19156 13376
rect 18380 13336 18386 13348
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 16945 13311 17003 13317
rect 16945 13308 16957 13311
rect 16592 13280 16957 13308
rect 16485 13271 16543 13277
rect 16945 13277 16957 13280
rect 16991 13277 17003 13311
rect 16945 13271 17003 13277
rect 17034 13268 17040 13320
rect 17092 13308 17098 13320
rect 17129 13311 17187 13317
rect 17129 13308 17141 13311
rect 17092 13280 17141 13308
rect 17092 13268 17098 13280
rect 17129 13277 17141 13280
rect 17175 13277 17187 13311
rect 17129 13271 17187 13277
rect 18046 13268 18052 13320
rect 18104 13308 18110 13320
rect 19812 13308 19840 13407
rect 20806 13404 20812 13416
rect 20864 13404 20870 13456
rect 21545 13447 21603 13453
rect 21545 13413 21557 13447
rect 21591 13444 21603 13447
rect 22094 13444 22100 13456
rect 21591 13416 22100 13444
rect 21591 13413 21603 13416
rect 21545 13407 21603 13413
rect 22094 13404 22100 13416
rect 22152 13404 22158 13456
rect 22480 13453 22508 13484
rect 22465 13447 22523 13453
rect 22465 13413 22477 13447
rect 22511 13413 22523 13447
rect 22465 13407 22523 13413
rect 20349 13379 20407 13385
rect 20349 13345 20361 13379
rect 20395 13376 20407 13379
rect 21358 13376 21364 13388
rect 20395 13348 21364 13376
rect 20395 13345 20407 13348
rect 20349 13339 20407 13345
rect 21358 13336 21364 13348
rect 21416 13336 21422 13388
rect 21634 13336 21640 13388
rect 21692 13376 21698 13388
rect 21729 13379 21787 13385
rect 21729 13376 21741 13379
rect 21692 13348 21741 13376
rect 21692 13336 21698 13348
rect 21729 13345 21741 13348
rect 21775 13376 21787 13379
rect 22002 13376 22008 13388
rect 21775 13348 22008 13376
rect 21775 13345 21787 13348
rect 21729 13339 21787 13345
rect 22002 13336 22008 13348
rect 22060 13336 22066 13388
rect 22112 13376 22140 13404
rect 22189 13379 22247 13385
rect 22189 13376 22201 13379
rect 22112 13348 22201 13376
rect 22189 13345 22201 13348
rect 22235 13345 22247 13379
rect 22189 13339 22247 13345
rect 22646 13336 22652 13388
rect 22704 13336 22710 13388
rect 18104 13280 19840 13308
rect 18104 13268 18110 13280
rect 20438 13268 20444 13320
rect 20496 13268 20502 13320
rect 20530 13268 20536 13320
rect 20588 13268 20594 13320
rect 20622 13268 20628 13320
rect 20680 13268 20686 13320
rect 17052 13240 17080 13268
rect 16592 13212 17080 13240
rect 18601 13243 18659 13249
rect 4890 13132 4896 13184
rect 4948 13132 4954 13184
rect 5810 13132 5816 13184
rect 5868 13132 5874 13184
rect 8113 13175 8171 13181
rect 8113 13141 8125 13175
rect 8159 13172 8171 13175
rect 8202 13172 8208 13184
rect 8159 13144 8208 13172
rect 8159 13141 8171 13144
rect 8113 13135 8171 13141
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 9122 13132 9128 13184
rect 9180 13132 9186 13184
rect 9306 13132 9312 13184
rect 9364 13132 9370 13184
rect 9766 13132 9772 13184
rect 9824 13132 9830 13184
rect 13541 13175 13599 13181
rect 13541 13141 13553 13175
rect 13587 13172 13599 13175
rect 13630 13172 13636 13184
rect 13587 13144 13636 13172
rect 13587 13141 13599 13144
rect 13541 13135 13599 13141
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 16592 13181 16620 13212
rect 18601 13209 18613 13243
rect 18647 13240 18659 13243
rect 19334 13240 19340 13252
rect 18647 13212 19340 13240
rect 18647 13209 18659 13212
rect 18601 13203 18659 13209
rect 19334 13200 19340 13212
rect 19392 13240 19398 13252
rect 20165 13243 20223 13249
rect 19392 13212 19932 13240
rect 19392 13200 19398 13212
rect 16577 13175 16635 13181
rect 16577 13141 16589 13175
rect 16623 13141 16635 13175
rect 16577 13135 16635 13141
rect 18417 13175 18475 13181
rect 18417 13141 18429 13175
rect 18463 13172 18475 13175
rect 18506 13172 18512 13184
rect 18463 13144 18512 13172
rect 18463 13141 18475 13144
rect 18417 13135 18475 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 19613 13175 19671 13181
rect 19613 13141 19625 13175
rect 19659 13172 19671 13175
rect 19702 13172 19708 13184
rect 19659 13144 19708 13172
rect 19659 13141 19671 13144
rect 19613 13135 19671 13141
rect 19702 13132 19708 13144
rect 19760 13132 19766 13184
rect 19794 13132 19800 13184
rect 19852 13132 19858 13184
rect 19904 13172 19932 13212
rect 20165 13209 20177 13243
rect 20211 13240 20223 13243
rect 20990 13240 20996 13252
rect 20211 13212 20996 13240
rect 20211 13209 20223 13212
rect 20165 13203 20223 13209
rect 20990 13200 20996 13212
rect 21048 13200 21054 13252
rect 21266 13200 21272 13252
rect 21324 13240 21330 13252
rect 22833 13243 22891 13249
rect 22833 13240 22845 13243
rect 21324 13212 22845 13240
rect 21324 13200 21330 13212
rect 22833 13209 22845 13212
rect 22879 13209 22891 13243
rect 22833 13203 22891 13209
rect 20622 13172 20628 13184
rect 19904 13144 20628 13172
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 20809 13175 20867 13181
rect 20809 13141 20821 13175
rect 20855 13172 20867 13175
rect 21082 13172 21088 13184
rect 20855 13144 21088 13172
rect 20855 13141 20867 13144
rect 20809 13135 20867 13141
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 21910 13132 21916 13184
rect 21968 13132 21974 13184
rect 552 13082 23368 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 23368 13082
rect 552 13008 23368 13030
rect 5902 12928 5908 12980
rect 5960 12968 5966 12980
rect 6178 12968 6184 12980
rect 5960 12940 6184 12968
rect 5960 12928 5966 12940
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 12342 12968 12348 12980
rect 11112 12940 12348 12968
rect 11112 12928 11118 12940
rect 8665 12835 8723 12841
rect 8665 12801 8677 12835
rect 8711 12832 8723 12835
rect 9030 12832 9036 12844
rect 8711 12804 9036 12832
rect 8711 12801 8723 12804
rect 8665 12795 8723 12801
rect 9030 12792 9036 12804
rect 9088 12832 9094 12844
rect 9217 12835 9275 12841
rect 9217 12832 9229 12835
rect 9088 12804 9229 12832
rect 9088 12792 9094 12804
rect 9217 12801 9229 12804
rect 9263 12801 9275 12835
rect 9217 12795 9275 12801
rect 11146 12792 11152 12844
rect 11204 12792 11210 12844
rect 11256 12841 11284 12940
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 12434 12928 12440 12980
rect 12492 12928 12498 12980
rect 15194 12968 15200 12980
rect 13556 12940 15200 12968
rect 13556 12900 13584 12940
rect 15194 12928 15200 12940
rect 15252 12928 15258 12980
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18693 12971 18751 12977
rect 18693 12968 18705 12971
rect 18095 12940 18705 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18693 12937 18705 12940
rect 18739 12937 18751 12971
rect 18693 12931 18751 12937
rect 20438 12928 20444 12980
rect 20496 12968 20502 12980
rect 20809 12971 20867 12977
rect 20809 12968 20821 12971
rect 20496 12940 20821 12968
rect 20496 12928 20502 12940
rect 20809 12937 20821 12940
rect 20855 12937 20867 12971
rect 20809 12931 20867 12937
rect 20898 12928 20904 12980
rect 20956 12928 20962 12980
rect 21082 12928 21088 12980
rect 21140 12928 21146 12980
rect 21358 12928 21364 12980
rect 21416 12968 21422 12980
rect 21729 12971 21787 12977
rect 21729 12968 21741 12971
rect 21416 12940 21741 12968
rect 21416 12928 21422 12940
rect 21729 12937 21741 12940
rect 21775 12937 21787 12971
rect 21729 12931 21787 12937
rect 11348 12872 13584 12900
rect 11241 12835 11299 12841
rect 11241 12801 11253 12835
rect 11287 12801 11299 12835
rect 11241 12795 11299 12801
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12733 4583 12767
rect 4525 12727 4583 12733
rect 4792 12767 4850 12773
rect 4792 12733 4804 12767
rect 4838 12764 4850 12767
rect 5810 12764 5816 12776
rect 4838 12736 5816 12764
rect 4838 12733 4850 12736
rect 4792 12727 4850 12733
rect 4246 12656 4252 12708
rect 4304 12696 4310 12708
rect 4540 12696 4568 12727
rect 5810 12724 5816 12736
rect 5868 12724 5874 12776
rect 5997 12767 6055 12773
rect 5997 12733 6009 12767
rect 6043 12733 6055 12767
rect 5997 12727 6055 12733
rect 5442 12696 5448 12708
rect 4304 12668 5448 12696
rect 4304 12656 4310 12668
rect 5442 12656 5448 12668
rect 5500 12696 5506 12708
rect 6012 12696 6040 12727
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 8444 12736 8585 12764
rect 8444 12724 8450 12736
rect 8573 12733 8585 12736
rect 8619 12733 8631 12767
rect 8573 12727 8631 12733
rect 8849 12767 8907 12773
rect 8849 12733 8861 12767
rect 8895 12764 8907 12767
rect 9122 12764 9128 12776
rect 8895 12736 9128 12764
rect 8895 12733 8907 12736
rect 8849 12727 8907 12733
rect 9122 12724 9128 12736
rect 9180 12724 9186 12776
rect 9306 12724 9312 12776
rect 9364 12724 9370 12776
rect 11348 12773 11376 12872
rect 18414 12860 18420 12912
rect 18472 12860 18478 12912
rect 21453 12903 21511 12909
rect 21453 12869 21465 12903
rect 21499 12900 21511 12903
rect 21913 12903 21971 12909
rect 21913 12900 21925 12903
rect 21499 12872 21925 12900
rect 21499 12869 21511 12872
rect 21453 12863 21511 12869
rect 18432 12832 18460 12860
rect 18432 12804 19196 12832
rect 11333 12767 11391 12773
rect 11333 12764 11345 12767
rect 10796 12736 11345 12764
rect 5500 12668 6040 12696
rect 6264 12699 6322 12705
rect 5500 12656 5506 12668
rect 6264 12665 6276 12699
rect 6310 12696 6322 12699
rect 6454 12696 6460 12708
rect 6310 12668 6460 12696
rect 6310 12665 6322 12668
rect 6264 12659 6322 12665
rect 6454 12656 6460 12668
rect 6512 12656 6518 12708
rect 6822 12656 6828 12708
rect 6880 12696 6886 12708
rect 9033 12699 9091 12705
rect 6880 12668 8984 12696
rect 6880 12656 6886 12668
rect 7374 12588 7380 12640
rect 7432 12588 7438 12640
rect 8956 12628 8984 12668
rect 9033 12665 9045 12699
rect 9079 12696 9091 12699
rect 9674 12696 9680 12708
rect 9079 12668 9680 12696
rect 9079 12665 9091 12668
rect 9033 12659 9091 12665
rect 9674 12656 9680 12668
rect 9732 12656 9738 12708
rect 10796 12640 10824 12736
rect 11333 12733 11345 12736
rect 11379 12733 11391 12767
rect 11333 12727 11391 12733
rect 11422 12724 11428 12776
rect 11480 12724 11486 12776
rect 11974 12724 11980 12776
rect 12032 12724 12038 12776
rect 12526 12724 12532 12776
rect 12584 12724 12590 12776
rect 13538 12724 13544 12776
rect 13596 12724 13602 12776
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 13797 12767 13855 12773
rect 13797 12764 13809 12767
rect 13688 12736 13809 12764
rect 13688 12724 13694 12736
rect 13797 12733 13809 12736
rect 13843 12733 13855 12767
rect 13797 12727 13855 12733
rect 18417 12767 18475 12773
rect 18417 12733 18429 12767
rect 18463 12733 18475 12767
rect 18417 12727 18475 12733
rect 11514 12656 11520 12708
rect 11572 12696 11578 12708
rect 12069 12699 12127 12705
rect 12069 12696 12081 12699
rect 11572 12668 12081 12696
rect 11572 12656 11578 12668
rect 12069 12665 12081 12668
rect 12115 12696 12127 12699
rect 12894 12696 12900 12708
rect 12115 12668 12900 12696
rect 12115 12665 12127 12668
rect 12069 12659 12127 12665
rect 12894 12656 12900 12668
rect 12952 12656 12958 12708
rect 18046 12656 18052 12708
rect 18104 12656 18110 12708
rect 18432 12696 18460 12727
rect 18506 12724 18512 12776
rect 18564 12764 18570 12776
rect 18877 12767 18935 12773
rect 18877 12764 18889 12767
rect 18564 12736 18889 12764
rect 18564 12724 18570 12736
rect 18877 12733 18889 12736
rect 18923 12764 18935 12767
rect 19058 12764 19064 12776
rect 18923 12736 19064 12764
rect 18923 12733 18935 12736
rect 18877 12727 18935 12733
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 19168 12773 19196 12804
rect 19153 12767 19211 12773
rect 19153 12733 19165 12767
rect 19199 12733 19211 12767
rect 19153 12727 19211 12733
rect 19426 12724 19432 12776
rect 19484 12724 19490 12776
rect 19702 12773 19708 12776
rect 19696 12764 19708 12773
rect 19663 12736 19708 12764
rect 19696 12727 19708 12736
rect 19702 12724 19708 12727
rect 19760 12724 19766 12776
rect 20714 12724 20720 12776
rect 20772 12764 20778 12776
rect 20772 12736 21588 12764
rect 20772 12724 20778 12736
rect 19334 12696 19340 12708
rect 18432 12668 19340 12696
rect 19334 12656 19340 12668
rect 19392 12656 19398 12708
rect 20990 12656 20996 12708
rect 21048 12696 21054 12708
rect 21560 12705 21588 12736
rect 21545 12699 21603 12705
rect 21048 12668 21220 12696
rect 21048 12656 21054 12668
rect 10778 12628 10784 12640
rect 8956 12600 10784 12628
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 10962 12588 10968 12640
rect 11020 12588 11026 12640
rect 12250 12588 12256 12640
rect 12308 12588 12314 12640
rect 14918 12588 14924 12640
rect 14976 12588 14982 12640
rect 17865 12631 17923 12637
rect 17865 12597 17877 12631
rect 17911 12628 17923 12631
rect 17954 12628 17960 12640
rect 17911 12600 17960 12628
rect 17911 12597 17923 12600
rect 17865 12591 17923 12597
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 19061 12631 19119 12637
rect 19061 12597 19073 12631
rect 19107 12628 19119 12631
rect 19150 12628 19156 12640
rect 19107 12600 19156 12628
rect 19107 12597 19119 12600
rect 19061 12591 19119 12597
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 21085 12631 21143 12637
rect 21085 12628 21097 12631
rect 20864 12600 21097 12628
rect 20864 12588 20870 12600
rect 21085 12597 21097 12600
rect 21131 12597 21143 12631
rect 21192 12628 21220 12668
rect 21545 12665 21557 12699
rect 21591 12665 21603 12699
rect 21744 12696 21772 12872
rect 21913 12869 21925 12872
rect 21959 12869 21971 12903
rect 21913 12863 21971 12869
rect 21818 12792 21824 12844
rect 21876 12832 21882 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21876 12804 22017 12832
rect 21876 12792 21882 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 22278 12724 22284 12776
rect 22336 12724 22342 12776
rect 22094 12696 22100 12708
rect 21744 12668 22100 12696
rect 21545 12659 21603 12665
rect 22094 12656 22100 12668
rect 22152 12656 22158 12708
rect 21745 12631 21803 12637
rect 21745 12628 21757 12631
rect 21192 12600 21757 12628
rect 21085 12591 21143 12597
rect 21745 12597 21757 12600
rect 21791 12597 21803 12631
rect 21745 12591 21803 12597
rect 552 12538 23368 12560
rect 552 12486 4322 12538
rect 4374 12486 4386 12538
rect 4438 12486 4450 12538
rect 4502 12486 4514 12538
rect 4566 12486 4578 12538
rect 4630 12486 23368 12538
rect 552 12464 23368 12486
rect 5258 12384 5264 12436
rect 5316 12424 5322 12436
rect 5629 12427 5687 12433
rect 5629 12424 5641 12427
rect 5316 12396 5641 12424
rect 5316 12384 5322 12396
rect 5629 12393 5641 12396
rect 5675 12393 5687 12427
rect 5629 12387 5687 12393
rect 6454 12384 6460 12436
rect 6512 12384 6518 12436
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 6696 12396 6929 12424
rect 6696 12384 6702 12396
rect 6917 12393 6929 12396
rect 6963 12393 6975 12427
rect 6917 12387 6975 12393
rect 11333 12427 11391 12433
rect 11333 12393 11345 12427
rect 11379 12424 11391 12427
rect 11422 12424 11428 12436
rect 11379 12396 11428 12424
rect 11379 12393 11391 12396
rect 11333 12387 11391 12393
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 13173 12427 13231 12433
rect 13173 12424 13185 12427
rect 12032 12396 13185 12424
rect 12032 12384 12038 12396
rect 13173 12393 13185 12396
rect 13219 12393 13231 12427
rect 13173 12387 13231 12393
rect 13998 12384 14004 12436
rect 14056 12424 14062 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 14056 12396 14105 12424
rect 14056 12384 14062 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 14093 12387 14151 12393
rect 14642 12384 14648 12436
rect 14700 12424 14706 12436
rect 15197 12427 15255 12433
rect 15197 12424 15209 12427
rect 14700 12396 15209 12424
rect 14700 12384 14706 12396
rect 15197 12393 15209 12396
rect 15243 12393 15255 12427
rect 15197 12387 15255 12393
rect 17589 12427 17647 12433
rect 17589 12393 17601 12427
rect 17635 12424 17647 12427
rect 17635 12396 18552 12424
rect 17635 12393 17647 12396
rect 17589 12387 17647 12393
rect 4516 12359 4574 12365
rect 4516 12325 4528 12359
rect 4562 12356 4574 12359
rect 4890 12356 4896 12368
rect 4562 12328 4896 12356
rect 4562 12325 4574 12328
rect 4516 12319 4574 12325
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 6825 12359 6883 12365
rect 6825 12325 6837 12359
rect 6871 12356 6883 12359
rect 7374 12356 7380 12368
rect 6871 12328 7380 12356
rect 6871 12325 6883 12328
rect 6825 12319 6883 12325
rect 7374 12316 7380 12328
rect 7432 12356 7438 12368
rect 7926 12356 7932 12368
rect 7432 12328 7932 12356
rect 7432 12316 7438 12328
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 8021 12359 8079 12365
rect 8021 12325 8033 12359
rect 8067 12356 8079 12359
rect 8386 12356 8392 12368
rect 8067 12328 8392 12356
rect 8067 12325 8079 12328
rect 8021 12319 8079 12325
rect 8386 12316 8392 12328
rect 8444 12316 8450 12368
rect 12060 12359 12118 12365
rect 8588 12328 11468 12356
rect 8588 12300 8616 12328
rect 4246 12248 4252 12300
rect 4304 12248 4310 12300
rect 8113 12291 8171 12297
rect 8113 12257 8125 12291
rect 8159 12257 8171 12291
rect 8113 12251 8171 12257
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12189 7067 12223
rect 8128 12220 8156 12251
rect 8202 12248 8208 12300
rect 8260 12248 8266 12300
rect 8478 12248 8484 12300
rect 8536 12248 8542 12300
rect 8570 12248 8576 12300
rect 8628 12248 8634 12300
rect 9214 12288 9220 12300
rect 8864 12260 9220 12288
rect 8864 12220 8892 12260
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 9766 12248 9772 12300
rect 9824 12248 9830 12300
rect 11440 12288 11468 12328
rect 12060 12325 12072 12359
rect 12106 12356 12118 12359
rect 12250 12356 12256 12368
rect 12106 12328 12256 12356
rect 12106 12325 12118 12328
rect 12060 12319 12118 12325
rect 12250 12316 12256 12328
rect 12308 12316 12314 12368
rect 16206 12356 16212 12368
rect 14292 12328 16212 12356
rect 11514 12288 11520 12300
rect 11440 12260 11520 12288
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 14292 12297 14320 12328
rect 16206 12316 16212 12328
rect 16264 12316 16270 12368
rect 17221 12359 17279 12365
rect 17221 12325 17233 12359
rect 17267 12356 17279 12359
rect 17310 12356 17316 12368
rect 17267 12328 17316 12356
rect 17267 12325 17279 12328
rect 17221 12319 17279 12325
rect 17310 12316 17316 12328
rect 17368 12316 17374 12368
rect 17437 12359 17495 12365
rect 17437 12325 17449 12359
rect 17483 12356 17495 12359
rect 17770 12356 17776 12368
rect 17483 12328 17776 12356
rect 17483 12325 17495 12328
rect 17437 12319 17495 12325
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 17954 12365 17960 12368
rect 17948 12356 17960 12365
rect 17915 12328 17960 12356
rect 17948 12319 17960 12328
rect 17954 12316 17960 12319
rect 18012 12316 18018 12368
rect 18046 12316 18052 12368
rect 18104 12316 18110 12368
rect 18524 12356 18552 12396
rect 19058 12384 19064 12436
rect 19116 12384 19122 12436
rect 19150 12384 19156 12436
rect 19208 12424 19214 12436
rect 20533 12427 20591 12433
rect 20533 12424 20545 12427
rect 19208 12396 20545 12424
rect 19208 12384 19214 12396
rect 20533 12393 20545 12396
rect 20579 12393 20591 12427
rect 20533 12387 20591 12393
rect 20990 12384 20996 12436
rect 21048 12384 21054 12436
rect 21634 12384 21640 12436
rect 21692 12384 21698 12436
rect 19398 12359 19456 12365
rect 19398 12356 19410 12359
rect 18524 12328 19410 12356
rect 19398 12325 19410 12328
rect 19444 12325 19456 12359
rect 19398 12319 19456 12325
rect 20622 12316 20628 12368
rect 20680 12316 20686 12368
rect 21358 12316 21364 12368
rect 21416 12356 21422 12368
rect 22278 12356 22284 12368
rect 21416 12328 22284 12356
rect 21416 12316 21422 12328
rect 22278 12316 22284 12328
rect 22336 12316 22342 12368
rect 11793 12291 11851 12297
rect 11793 12288 11805 12291
rect 11624 12260 11805 12288
rect 8128 12192 8892 12220
rect 7009 12183 7067 12189
rect 6822 12112 6828 12164
rect 6880 12152 6886 12164
rect 7024 12152 7052 12183
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 9088 12192 9137 12220
rect 9088 12180 9094 12192
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9674 12180 9680 12232
rect 9732 12180 9738 12232
rect 10686 12180 10692 12232
rect 10744 12220 10750 12232
rect 11624 12220 11652 12260
rect 11793 12257 11805 12260
rect 11839 12257 11851 12291
rect 11793 12251 11851 12257
rect 14277 12291 14335 12297
rect 14277 12257 14289 12291
rect 14323 12257 14335 12291
rect 14277 12251 14335 12257
rect 14461 12291 14519 12297
rect 14461 12257 14473 12291
rect 14507 12288 14519 12291
rect 14918 12288 14924 12300
rect 14507 12260 14924 12288
rect 14507 12257 14519 12260
rect 14461 12251 14519 12257
rect 14918 12248 14924 12260
rect 14976 12248 14982 12300
rect 15102 12248 15108 12300
rect 15160 12248 15166 12300
rect 16298 12248 16304 12300
rect 16356 12248 16362 12300
rect 16942 12248 16948 12300
rect 17000 12248 17006 12300
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12288 17187 12291
rect 18064 12288 18092 12316
rect 17175 12260 18092 12288
rect 17175 12257 17187 12260
rect 17129 12251 17187 12257
rect 20254 12248 20260 12300
rect 20312 12288 20318 12300
rect 20640 12288 20668 12316
rect 20809 12291 20867 12297
rect 20809 12288 20821 12291
rect 20312 12260 20821 12288
rect 20312 12248 20318 12260
rect 20809 12257 20821 12260
rect 20855 12257 20867 12291
rect 20809 12251 20867 12257
rect 22002 12248 22008 12300
rect 22060 12288 22066 12300
rect 22750 12291 22808 12297
rect 22750 12288 22762 12291
rect 22060 12260 22762 12288
rect 22060 12248 22066 12260
rect 22750 12257 22762 12260
rect 22796 12257 22808 12291
rect 22750 12251 22808 12257
rect 10744 12192 11652 12220
rect 10744 12180 10750 12192
rect 11698 12180 11704 12232
rect 11756 12180 11762 12232
rect 14550 12180 14556 12232
rect 14608 12220 14614 12232
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 14608 12192 15301 12220
rect 14608 12180 14614 12192
rect 15289 12189 15301 12192
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 16390 12180 16396 12232
rect 16448 12180 16454 12232
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12189 17739 12223
rect 17681 12183 17739 12189
rect 6880 12124 7052 12152
rect 10137 12155 10195 12161
rect 6880 12112 6886 12124
rect 10137 12121 10149 12155
rect 10183 12152 10195 12155
rect 10870 12152 10876 12164
rect 10183 12124 10876 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 10870 12112 10876 12124
rect 10928 12112 10934 12164
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 8757 12087 8815 12093
rect 8757 12084 8769 12087
rect 8720 12056 8769 12084
rect 8720 12044 8726 12056
rect 8757 12053 8769 12056
rect 8803 12053 8815 12087
rect 8757 12047 8815 12053
rect 8938 12044 8944 12096
rect 8996 12044 9002 12096
rect 14642 12044 14648 12096
rect 14700 12084 14706 12096
rect 14737 12087 14795 12093
rect 14737 12084 14749 12087
rect 14700 12056 14749 12084
rect 14700 12044 14706 12056
rect 14737 12053 14749 12056
rect 14783 12053 14795 12087
rect 14737 12047 14795 12053
rect 16666 12044 16672 12096
rect 16724 12044 16730 12096
rect 17037 12087 17095 12093
rect 17037 12053 17049 12087
rect 17083 12084 17095 12087
rect 17405 12087 17463 12093
rect 17405 12084 17417 12087
rect 17083 12056 17417 12084
rect 17083 12053 17095 12056
rect 17037 12047 17095 12053
rect 17405 12053 17417 12056
rect 17451 12053 17463 12087
rect 17696 12084 17724 12183
rect 18690 12180 18696 12232
rect 18748 12220 18754 12232
rect 19153 12223 19211 12229
rect 19153 12220 19165 12223
rect 18748 12192 19165 12220
rect 18748 12180 18754 12192
rect 19153 12189 19165 12192
rect 19199 12189 19211 12223
rect 19153 12183 19211 12189
rect 20438 12180 20444 12232
rect 20496 12220 20502 12232
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 20496 12192 20637 12220
rect 20496 12180 20502 12192
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 23017 12223 23075 12229
rect 23017 12189 23029 12223
rect 23063 12220 23075 12223
rect 23063 12192 23428 12220
rect 23063 12189 23075 12192
rect 23017 12183 23075 12189
rect 19426 12084 19432 12096
rect 17696 12056 19432 12084
rect 17405 12047 17463 12053
rect 19426 12044 19432 12056
rect 19484 12044 19490 12096
rect 20162 12044 20168 12096
rect 20220 12084 20226 12096
rect 21453 12087 21511 12093
rect 21453 12084 21465 12087
rect 20220 12056 21465 12084
rect 20220 12044 20226 12056
rect 21453 12053 21465 12056
rect 21499 12053 21511 12087
rect 21453 12047 21511 12053
rect 552 11994 23368 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 23368 11994
rect 552 11920 23368 11942
rect 5626 11840 5632 11892
rect 5684 11840 5690 11892
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 9582 11880 9588 11892
rect 8628 11852 9588 11880
rect 8628 11840 8634 11852
rect 9582 11840 9588 11852
rect 9640 11880 9646 11892
rect 9769 11883 9827 11889
rect 9769 11880 9781 11883
rect 9640 11852 9781 11880
rect 9640 11840 9646 11852
rect 9769 11849 9781 11852
rect 9815 11849 9827 11883
rect 9769 11843 9827 11849
rect 11698 11840 11704 11892
rect 11756 11880 11762 11892
rect 12066 11880 12072 11892
rect 11756 11852 12072 11880
rect 11756 11840 11762 11852
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 14185 11883 14243 11889
rect 14185 11849 14197 11883
rect 14231 11880 14243 11883
rect 14550 11880 14556 11892
rect 14231 11852 14556 11880
rect 14231 11849 14243 11852
rect 14185 11843 14243 11849
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 15102 11840 15108 11892
rect 15160 11880 15166 11892
rect 15749 11883 15807 11889
rect 15749 11880 15761 11883
rect 15160 11852 15761 11880
rect 15160 11840 15166 11852
rect 15749 11849 15761 11852
rect 15795 11849 15807 11883
rect 15749 11843 15807 11849
rect 17770 11840 17776 11892
rect 17828 11880 17834 11892
rect 17865 11883 17923 11889
rect 17865 11880 17877 11883
rect 17828 11852 17877 11880
rect 17828 11840 17834 11852
rect 17865 11849 17877 11852
rect 17911 11849 17923 11883
rect 17865 11843 17923 11849
rect 19705 11883 19763 11889
rect 19705 11849 19717 11883
rect 19751 11880 19763 11883
rect 19794 11880 19800 11892
rect 19751 11852 19800 11880
rect 19751 11849 19763 11852
rect 19705 11843 19763 11849
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 21266 11840 21272 11892
rect 21324 11840 21330 11892
rect 23400 11880 23428 12192
rect 21560 11852 23428 11880
rect 5534 11772 5540 11824
rect 5592 11772 5598 11824
rect 19426 11772 19432 11824
rect 19484 11812 19490 11824
rect 21560 11812 21588 11852
rect 19484 11784 21588 11812
rect 19484 11772 19490 11784
rect 5258 11704 5264 11756
rect 5316 11744 5322 11756
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5316 11716 5457 11744
rect 5316 11704 5322 11716
rect 5445 11713 5457 11716
rect 5491 11744 5503 11747
rect 5994 11744 6000 11756
rect 5491 11716 6000 11744
rect 5491 11713 5503 11716
rect 5445 11707 5503 11713
rect 5994 11704 6000 11716
rect 6052 11704 6058 11756
rect 20990 11744 20996 11756
rect 20548 11716 20996 11744
rect 5166 11636 5172 11688
rect 5224 11676 5230 11688
rect 5721 11679 5779 11685
rect 5721 11676 5733 11679
rect 5224 11648 5733 11676
rect 5224 11636 5230 11648
rect 5721 11645 5733 11648
rect 5767 11645 5779 11679
rect 5721 11639 5779 11645
rect 8386 11636 8392 11688
rect 8444 11636 8450 11688
rect 8662 11685 8668 11688
rect 8656 11676 8668 11685
rect 8623 11648 8668 11676
rect 8656 11639 8668 11648
rect 8662 11636 8668 11639
rect 8720 11636 8726 11688
rect 10686 11636 10692 11688
rect 10744 11636 10750 11688
rect 10962 11685 10968 11688
rect 10956 11639 10968 11685
rect 10962 11636 10968 11639
rect 11020 11636 11026 11688
rect 14001 11679 14059 11685
rect 14001 11645 14013 11679
rect 14047 11676 14059 11679
rect 14090 11676 14096 11688
rect 14047 11648 14096 11676
rect 14047 11645 14059 11648
rect 14001 11639 14059 11645
rect 14090 11636 14096 11648
rect 14148 11636 14154 11688
rect 14274 11636 14280 11688
rect 14332 11636 14338 11688
rect 14642 11685 14648 11688
rect 14369 11679 14427 11685
rect 14369 11645 14381 11679
rect 14415 11645 14427 11679
rect 14636 11676 14648 11685
rect 14603 11648 14648 11676
rect 14369 11639 14427 11645
rect 14636 11639 14648 11648
rect 13446 11568 13452 11620
rect 13504 11608 13510 11620
rect 14384 11608 14412 11639
rect 14642 11636 14648 11639
rect 14700 11636 14706 11688
rect 18046 11636 18052 11688
rect 18104 11676 18110 11688
rect 19150 11676 19156 11688
rect 18104 11648 19156 11676
rect 18104 11636 18110 11648
rect 19150 11636 19156 11648
rect 19208 11636 19214 11688
rect 19889 11679 19947 11685
rect 19889 11645 19901 11679
rect 19935 11676 19947 11679
rect 20438 11676 20444 11688
rect 19935 11648 20444 11676
rect 19935 11645 19947 11648
rect 19889 11639 19947 11645
rect 20438 11636 20444 11648
rect 20496 11636 20502 11688
rect 20548 11685 20576 11716
rect 20533 11679 20591 11685
rect 20533 11645 20545 11679
rect 20579 11645 20591 11679
rect 20533 11639 20591 11645
rect 20625 11679 20683 11685
rect 20625 11645 20637 11679
rect 20671 11676 20683 11679
rect 20714 11676 20720 11688
rect 20671 11648 20720 11676
rect 20671 11645 20683 11648
rect 20625 11639 20683 11645
rect 15010 11608 15016 11620
rect 13504 11580 15016 11608
rect 13504 11568 13510 11580
rect 15010 11568 15016 11580
rect 15068 11568 15074 11620
rect 18233 11611 18291 11617
rect 18233 11577 18245 11611
rect 18279 11608 18291 11611
rect 18414 11608 18420 11620
rect 18279 11580 18420 11608
rect 18279 11577 18291 11580
rect 18233 11571 18291 11577
rect 18414 11568 18420 11580
rect 18472 11568 18478 11620
rect 20073 11611 20131 11617
rect 20073 11577 20085 11611
rect 20119 11608 20131 11611
rect 20254 11608 20260 11620
rect 20119 11580 20260 11608
rect 20119 11577 20131 11580
rect 20073 11571 20131 11577
rect 20254 11568 20260 11580
rect 20312 11568 20318 11620
rect 20349 11611 20407 11617
rect 20349 11577 20361 11611
rect 20395 11608 20407 11611
rect 20640 11608 20668 11639
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 20824 11685 20852 11716
rect 20990 11704 20996 11716
rect 21048 11704 21054 11756
rect 21560 11753 21588 11784
rect 21545 11747 21603 11753
rect 21545 11713 21557 11747
rect 21591 11713 21603 11747
rect 21545 11707 21603 11713
rect 20809 11679 20867 11685
rect 20809 11645 20821 11679
rect 20855 11645 20867 11679
rect 20809 11639 20867 11645
rect 20901 11679 20959 11685
rect 20901 11645 20913 11679
rect 20947 11676 20959 11679
rect 21082 11676 21088 11688
rect 20947 11648 21088 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 21082 11636 21088 11648
rect 21140 11636 21146 11688
rect 21790 11611 21848 11617
rect 21790 11608 21802 11611
rect 20395 11580 20668 11608
rect 21468 11580 21802 11608
rect 20395 11577 20407 11580
rect 20349 11571 20407 11577
rect 13814 11500 13820 11552
rect 13872 11500 13878 11552
rect 19978 11500 19984 11552
rect 20036 11540 20042 11552
rect 20165 11543 20223 11549
rect 20165 11540 20177 11543
rect 20036 11512 20177 11540
rect 20036 11500 20042 11512
rect 20165 11509 20177 11512
rect 20211 11509 20223 11543
rect 20165 11503 20223 11509
rect 20714 11500 20720 11552
rect 20772 11500 20778 11552
rect 20990 11500 20996 11552
rect 21048 11540 21054 11552
rect 21468 11549 21496 11580
rect 21790 11577 21802 11580
rect 21836 11577 21848 11611
rect 21790 11571 21848 11577
rect 21269 11543 21327 11549
rect 21269 11540 21281 11543
rect 21048 11512 21281 11540
rect 21048 11500 21054 11512
rect 21269 11509 21281 11512
rect 21315 11509 21327 11543
rect 21269 11503 21327 11509
rect 21453 11543 21511 11549
rect 21453 11509 21465 11543
rect 21499 11509 21511 11543
rect 21453 11503 21511 11509
rect 22278 11500 22284 11552
rect 22336 11540 22342 11552
rect 22646 11540 22652 11552
rect 22336 11512 22652 11540
rect 22336 11500 22342 11512
rect 22646 11500 22652 11512
rect 22704 11540 22710 11552
rect 22925 11543 22983 11549
rect 22925 11540 22937 11543
rect 22704 11512 22937 11540
rect 22704 11500 22710 11512
rect 22925 11509 22937 11512
rect 22971 11509 22983 11543
rect 22925 11503 22983 11509
rect 552 11450 23368 11472
rect 552 11398 4322 11450
rect 4374 11398 4386 11450
rect 4438 11398 4450 11450
rect 4502 11398 4514 11450
rect 4566 11398 4578 11450
rect 4630 11398 23368 11450
rect 552 11376 23368 11398
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 7837 11339 7895 11345
rect 7837 11336 7849 11339
rect 5500 11308 7849 11336
rect 5500 11296 5506 11308
rect 7837 11305 7849 11308
rect 7883 11336 7895 11339
rect 8386 11336 8392 11348
rect 7883 11308 8392 11336
rect 7883 11305 7895 11308
rect 7837 11299 7895 11305
rect 5166 11228 5172 11280
rect 5224 11228 5230 11280
rect 5902 11228 5908 11280
rect 5960 11268 5966 11280
rect 6270 11268 6276 11280
rect 5960 11240 6276 11268
rect 5960 11228 5966 11240
rect 6270 11228 6276 11240
rect 6328 11228 6334 11280
rect 8036 11268 8064 11308
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 14274 11296 14280 11348
rect 14332 11336 14338 11348
rect 14829 11339 14887 11345
rect 14829 11336 14841 11339
rect 14332 11308 14841 11336
rect 14332 11296 14338 11308
rect 14829 11305 14841 11308
rect 14875 11305 14887 11339
rect 14829 11299 14887 11305
rect 10686 11268 10692 11280
rect 8036 11240 8156 11268
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5184 11200 5212 11228
rect 8128 11209 8156 11240
rect 8220 11240 10692 11268
rect 6181 11203 6239 11209
rect 6181 11200 6193 11203
rect 5123 11172 6193 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 6181 11169 6193 11172
rect 6227 11169 6239 11203
rect 6181 11163 6239 11169
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 8113 11203 8171 11209
rect 8113 11169 8125 11203
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 5718 11132 5724 11144
rect 5215 11104 5724 11132
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 5718 11092 5724 11104
rect 5776 11092 5782 11144
rect 5994 11092 6000 11144
rect 6052 11092 6058 11144
rect 8036 11132 8064 11163
rect 8220 11132 8248 11240
rect 10686 11228 10692 11240
rect 10744 11268 10750 11280
rect 13716 11271 13774 11277
rect 10744 11240 11008 11268
rect 10744 11228 10750 11240
rect 10980 11212 11008 11240
rect 13716 11237 13728 11271
rect 13762 11268 13774 11271
rect 13814 11268 13820 11280
rect 13762 11240 13820 11268
rect 13762 11237 13774 11240
rect 13716 11231 13774 11237
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 8380 11203 8438 11209
rect 8380 11169 8392 11203
rect 8426 11200 8438 11203
rect 8662 11200 8668 11212
rect 8426 11172 8668 11200
rect 8426 11169 8438 11172
rect 8380 11163 8438 11169
rect 8662 11160 8668 11172
rect 8720 11160 8726 11212
rect 10962 11160 10968 11212
rect 11020 11160 11026 11212
rect 11238 11209 11244 11212
rect 11232 11163 11244 11209
rect 11238 11160 11244 11163
rect 11296 11160 11302 11212
rect 13446 11160 13452 11212
rect 13504 11160 13510 11212
rect 8036 11104 8248 11132
rect 5445 11067 5503 11073
rect 5445 11033 5457 11067
rect 5491 11064 5503 11067
rect 5626 11064 5632 11076
rect 5491 11036 5632 11064
rect 5491 11033 5503 11036
rect 5445 11027 5503 11033
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 6365 11067 6423 11073
rect 6365 11033 6377 11067
rect 6411 11064 6423 11067
rect 7006 11064 7012 11076
rect 6411 11036 7012 11064
rect 6411 11033 6423 11036
rect 6365 11027 6423 11033
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 5718 10956 5724 11008
rect 5776 10996 5782 11008
rect 5905 10999 5963 11005
rect 5905 10996 5917 10999
rect 5776 10968 5917 10996
rect 5776 10956 5782 10968
rect 5905 10965 5917 10968
rect 5951 10965 5963 10999
rect 5905 10959 5963 10965
rect 9490 10956 9496 11008
rect 9548 10956 9554 11008
rect 12342 10956 12348 11008
rect 12400 10956 12406 11008
rect 14844 10996 14872 11299
rect 14918 11296 14924 11348
rect 14976 11296 14982 11348
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 17865 11339 17923 11345
rect 17865 11336 17877 11339
rect 17368 11308 17877 11336
rect 17368 11296 17374 11308
rect 17865 11305 17877 11308
rect 17911 11336 17923 11339
rect 20162 11336 20168 11348
rect 17911 11308 20168 11336
rect 17911 11305 17923 11308
rect 17865 11299 17923 11305
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 20806 11296 20812 11348
rect 20864 11296 20870 11348
rect 21634 11296 21640 11348
rect 21692 11336 21698 11348
rect 21692 11308 21956 11336
rect 21692 11296 21698 11308
rect 14936 11268 14964 11296
rect 14936 11240 15240 11268
rect 14918 11160 14924 11212
rect 14976 11160 14982 11212
rect 15102 11160 15108 11212
rect 15160 11160 15166 11212
rect 15212 11209 15240 11240
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 17189 11271 17247 11277
rect 17189 11268 17201 11271
rect 16264 11240 17201 11268
rect 16264 11228 16270 11240
rect 17189 11237 17201 11240
rect 17235 11237 17247 11271
rect 17189 11231 17247 11237
rect 17405 11271 17463 11277
rect 17405 11237 17417 11271
rect 17451 11268 17463 11271
rect 17770 11268 17776 11280
rect 17451 11240 17776 11268
rect 17451 11237 17463 11240
rect 17405 11231 17463 11237
rect 17770 11228 17776 11240
rect 17828 11228 17834 11280
rect 20180 11268 20208 11296
rect 21821 11271 21879 11277
rect 21821 11268 21833 11271
rect 20180 11240 21833 11268
rect 21821 11237 21833 11240
rect 21867 11237 21879 11271
rect 21928 11268 21956 11308
rect 22002 11296 22008 11348
rect 22060 11296 22066 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 22255 11339 22313 11345
rect 22255 11336 22267 11339
rect 22152 11308 22267 11336
rect 22152 11296 22158 11308
rect 22255 11305 22267 11308
rect 22301 11305 22313 11339
rect 22255 11299 22313 11305
rect 22465 11271 22523 11277
rect 22465 11268 22477 11271
rect 21928 11240 22477 11268
rect 21821 11231 21879 11237
rect 22465 11237 22477 11240
rect 22511 11237 22523 11271
rect 22465 11231 22523 11237
rect 15197 11203 15255 11209
rect 15197 11169 15209 11203
rect 15243 11169 15255 11203
rect 15197 11163 15255 11169
rect 16574 11160 16580 11212
rect 16632 11160 16638 11212
rect 16942 11160 16948 11212
rect 17000 11200 17006 11212
rect 17497 11203 17555 11209
rect 17497 11200 17509 11203
rect 17000 11172 17509 11200
rect 17000 11160 17006 11172
rect 17497 11169 17509 11172
rect 17543 11200 17555 11203
rect 18414 11200 18420 11212
rect 17543 11172 18420 11200
rect 17543 11169 17555 11172
rect 17497 11163 17555 11169
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 19426 11160 19432 11212
rect 19484 11160 19490 11212
rect 19702 11209 19708 11212
rect 19696 11163 19708 11209
rect 19702 11160 19708 11163
rect 19760 11160 19766 11212
rect 21453 11203 21511 11209
rect 21453 11169 21465 11203
rect 21499 11200 21511 11203
rect 21726 11200 21732 11212
rect 21499 11172 21732 11200
rect 21499 11169 21511 11172
rect 21453 11163 21511 11169
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 21836 11200 21864 11231
rect 22741 11203 22799 11209
rect 22741 11200 22753 11203
rect 21836 11172 22753 11200
rect 22741 11169 22753 11172
rect 22787 11169 22799 11203
rect 22741 11163 22799 11169
rect 16666 11092 16672 11144
rect 16724 11092 16730 11144
rect 20990 11092 20996 11144
rect 21048 11132 21054 11144
rect 22557 11135 22615 11141
rect 22557 11132 22569 11135
rect 21048 11104 22569 11132
rect 21048 11092 21054 11104
rect 22557 11101 22569 11104
rect 22603 11101 22615 11135
rect 22557 11095 22615 11101
rect 15381 11067 15439 11073
rect 15381 11033 15393 11067
rect 15427 11064 15439 11067
rect 16390 11064 16396 11076
rect 15427 11036 16396 11064
rect 15427 11033 15439 11036
rect 15381 11027 15439 11033
rect 16390 11024 16396 11036
rect 16448 11064 16454 11076
rect 16448 11036 17172 11064
rect 16448 11024 16454 11036
rect 14921 10999 14979 11005
rect 14921 10996 14933 10999
rect 14844 10968 14933 10996
rect 14921 10965 14933 10968
rect 14967 10965 14979 10999
rect 14921 10959 14979 10965
rect 16850 10956 16856 11008
rect 16908 10956 16914 11008
rect 17034 10956 17040 11008
rect 17092 10956 17098 11008
rect 17144 10996 17172 11036
rect 20806 11024 20812 11076
rect 20864 11064 20870 11076
rect 21358 11064 21364 11076
rect 20864 11036 21364 11064
rect 20864 11024 20870 11036
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 17221 10999 17279 11005
rect 17221 10996 17233 10999
rect 17144 10968 17233 10996
rect 17221 10965 17233 10968
rect 17267 10965 17279 10999
rect 17221 10959 17279 10965
rect 17862 10956 17868 11008
rect 17920 10956 17926 11008
rect 18049 10999 18107 11005
rect 18049 10965 18061 10999
rect 18095 10996 18107 10999
rect 18230 10996 18236 11008
rect 18095 10968 18236 10996
rect 18095 10965 18107 10968
rect 18049 10959 18107 10965
rect 18230 10956 18236 10968
rect 18288 10956 18294 11008
rect 21821 10999 21879 11005
rect 21821 10965 21833 10999
rect 21867 10996 21879 10999
rect 21910 10996 21916 11008
rect 21867 10968 21916 10996
rect 21867 10965 21879 10968
rect 21821 10959 21879 10965
rect 21910 10956 21916 10968
rect 21968 10956 21974 11008
rect 22002 10956 22008 11008
rect 22060 10996 22066 11008
rect 22097 10999 22155 11005
rect 22097 10996 22109 10999
rect 22060 10968 22109 10996
rect 22060 10956 22066 10968
rect 22097 10965 22109 10968
rect 22143 10965 22155 10999
rect 22097 10959 22155 10965
rect 22278 10956 22284 11008
rect 22336 10956 22342 11008
rect 552 10906 23368 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 23368 10906
rect 552 10832 23368 10854
rect 5353 10795 5411 10801
rect 5353 10761 5365 10795
rect 5399 10792 5411 10795
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5399 10764 5641 10792
rect 5399 10761 5411 10764
rect 5353 10755 5411 10761
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 5629 10755 5687 10761
rect 5537 10727 5595 10733
rect 5537 10693 5549 10727
rect 5583 10693 5595 10727
rect 5644 10724 5672 10755
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 5813 10795 5871 10801
rect 5813 10792 5825 10795
rect 5776 10764 5825 10792
rect 5776 10752 5782 10764
rect 5813 10761 5825 10764
rect 5859 10761 5871 10795
rect 5813 10755 5871 10761
rect 6549 10795 6607 10801
rect 6549 10761 6561 10795
rect 6595 10792 6607 10795
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 6595 10764 7113 10792
rect 6595 10761 6607 10764
rect 6549 10755 6607 10761
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 7101 10755 7159 10761
rect 8662 10752 8668 10804
rect 8720 10752 8726 10804
rect 9582 10752 9588 10804
rect 9640 10752 9646 10804
rect 9953 10795 10011 10801
rect 9953 10761 9965 10795
rect 9999 10792 10011 10795
rect 9999 10764 11192 10792
rect 9999 10761 10011 10764
rect 9953 10755 10011 10761
rect 6733 10727 6791 10733
rect 5644 10696 6684 10724
rect 5537 10687 5595 10693
rect 5166 10616 5172 10668
rect 5224 10656 5230 10668
rect 5350 10656 5356 10668
rect 5224 10628 5356 10656
rect 5224 10616 5230 10628
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5552 10656 5580 10687
rect 6656 10656 6684 10696
rect 6733 10693 6745 10727
rect 6779 10724 6791 10727
rect 7190 10724 7196 10736
rect 6779 10696 7196 10724
rect 6779 10693 6791 10696
rect 6733 10687 6791 10693
rect 7190 10684 7196 10696
rect 7248 10684 7254 10736
rect 11164 10724 11192 10764
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11333 10795 11391 10801
rect 11333 10792 11345 10795
rect 11296 10764 11345 10792
rect 11296 10752 11302 10764
rect 11333 10761 11345 10764
rect 11379 10761 11391 10795
rect 11333 10755 11391 10761
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11655 10795 11713 10801
rect 11655 10792 11667 10795
rect 11480 10764 11667 10792
rect 11480 10752 11486 10764
rect 11655 10761 11667 10764
rect 11701 10792 11713 10795
rect 12066 10792 12072 10804
rect 11701 10764 12072 10792
rect 11701 10761 11713 10764
rect 11655 10755 11713 10761
rect 12066 10752 12072 10764
rect 12124 10752 12130 10804
rect 12529 10795 12587 10801
rect 12529 10761 12541 10795
rect 12575 10792 12587 10795
rect 12575 10764 13308 10792
rect 12575 10761 12587 10764
rect 12529 10755 12587 10761
rect 11793 10727 11851 10733
rect 11793 10724 11805 10727
rect 9324 10696 10824 10724
rect 11164 10696 11805 10724
rect 5552 10628 6592 10656
rect 6656 10628 6960 10656
rect 5184 10588 5212 10616
rect 5813 10591 5871 10597
rect 5813 10588 5825 10591
rect 5184 10560 5825 10588
rect 5813 10557 5825 10560
rect 5859 10557 5871 10591
rect 5813 10551 5871 10557
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 5997 10591 6055 10597
rect 5997 10588 6009 10591
rect 5960 10560 6009 10588
rect 5960 10548 5966 10560
rect 5997 10557 6009 10560
rect 6043 10557 6055 10591
rect 5997 10551 6055 10557
rect 6362 10548 6368 10600
rect 6420 10548 6426 10600
rect 6564 10597 6592 10628
rect 6932 10597 6960 10628
rect 8938 10616 8944 10668
rect 8996 10656 9002 10668
rect 9324 10665 9352 10696
rect 10796 10668 10824 10696
rect 11793 10693 11805 10696
rect 11839 10693 11851 10727
rect 11793 10687 11851 10693
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 8996 10628 9137 10656
rect 8996 10616 9002 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 9490 10616 9496 10668
rect 9548 10656 9554 10668
rect 9585 10659 9643 10665
rect 9585 10656 9597 10659
rect 9548 10628 9597 10656
rect 9548 10616 9554 10628
rect 9585 10625 9597 10628
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 10778 10616 10784 10668
rect 10836 10616 10842 10668
rect 10870 10616 10876 10668
rect 10928 10616 10934 10668
rect 6549 10591 6607 10597
rect 6549 10557 6561 10591
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10588 6975 10591
rect 7193 10591 7251 10597
rect 7193 10588 7205 10591
rect 6963 10560 7205 10588
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 7193 10557 7205 10560
rect 7239 10557 7251 10591
rect 7193 10551 7251 10557
rect 7377 10591 7435 10597
rect 7377 10557 7389 10591
rect 7423 10557 7435 10591
rect 7377 10551 7435 10557
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10588 9091 10591
rect 9508 10588 9536 10616
rect 9769 10591 9827 10597
rect 9769 10588 9781 10591
rect 9079 10560 9536 10588
rect 9600 10560 9781 10588
rect 9079 10557 9091 10560
rect 9033 10551 9091 10557
rect 5074 10480 5080 10532
rect 5132 10520 5138 10532
rect 5169 10523 5227 10529
rect 5169 10520 5181 10523
rect 5132 10492 5181 10520
rect 5132 10480 5138 10492
rect 5169 10489 5181 10492
rect 5215 10489 5227 10523
rect 5169 10483 5227 10489
rect 5385 10523 5443 10529
rect 5385 10489 5397 10523
rect 5431 10520 5443 10523
rect 5534 10520 5540 10532
rect 5431 10492 5540 10520
rect 5431 10489 5443 10492
rect 5385 10483 5443 10489
rect 5534 10480 5540 10492
rect 5592 10480 5598 10532
rect 6086 10480 6092 10532
rect 6144 10480 6150 10532
rect 6840 10520 6868 10551
rect 6196 10492 6868 10520
rect 5552 10452 5580 10480
rect 6196 10452 6224 10492
rect 7098 10480 7104 10532
rect 7156 10480 7162 10532
rect 7392 10520 7420 10551
rect 7208 10492 7420 10520
rect 5552 10424 6224 10452
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 7208 10452 7236 10492
rect 8938 10480 8944 10532
rect 8996 10520 9002 10532
rect 9493 10523 9551 10529
rect 9493 10520 9505 10523
rect 8996 10492 9505 10520
rect 8996 10480 9002 10492
rect 9493 10489 9505 10492
rect 9539 10489 9551 10523
rect 9493 10483 9551 10489
rect 6328 10424 7236 10452
rect 6328 10412 6334 10424
rect 7282 10412 7288 10464
rect 7340 10412 7346 10464
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 9600 10452 9628 10560
rect 9769 10557 9781 10560
rect 9815 10557 9827 10591
rect 9769 10551 9827 10557
rect 10965 10591 11023 10597
rect 10965 10557 10977 10591
rect 11011 10588 11023 10591
rect 11514 10588 11520 10600
rect 11011 10560 11520 10588
rect 11011 10557 11023 10560
rect 10965 10551 11023 10557
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 11808 10520 11836 10687
rect 12434 10684 12440 10736
rect 12492 10724 12498 10736
rect 12492 10696 13124 10724
rect 12492 10684 12498 10696
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 12268 10628 12756 10656
rect 11974 10548 11980 10600
rect 12032 10588 12038 10600
rect 12176 10588 12204 10619
rect 12032 10560 12204 10588
rect 12032 10548 12038 10560
rect 12066 10520 12072 10532
rect 11808 10492 12072 10520
rect 12066 10480 12072 10492
rect 12124 10520 12130 10532
rect 12268 10520 12296 10628
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 12728 10597 12756 10628
rect 13096 10597 13124 10696
rect 13280 10597 13308 10764
rect 14274 10752 14280 10804
rect 14332 10792 14338 10804
rect 14783 10795 14841 10801
rect 14783 10792 14795 10795
rect 14332 10764 14795 10792
rect 14332 10752 14338 10764
rect 14783 10761 14795 10764
rect 14829 10761 14841 10795
rect 14783 10755 14841 10761
rect 16853 10795 16911 10801
rect 16853 10761 16865 10795
rect 16899 10792 16911 10795
rect 17034 10792 17040 10804
rect 16899 10764 17040 10792
rect 16899 10761 16911 10764
rect 16853 10755 16911 10761
rect 17034 10752 17040 10764
rect 17092 10752 17098 10804
rect 17129 10795 17187 10801
rect 17129 10761 17141 10795
rect 17175 10792 17187 10795
rect 17218 10792 17224 10804
rect 17175 10764 17224 10792
rect 17175 10761 17187 10764
rect 17129 10755 17187 10761
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 19702 10752 19708 10804
rect 19760 10792 19766 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 19760 10764 19809 10792
rect 19760 10752 19766 10764
rect 19797 10761 19809 10764
rect 19843 10761 19855 10795
rect 19797 10755 19855 10761
rect 19981 10795 20039 10801
rect 19981 10761 19993 10795
rect 20027 10792 20039 10795
rect 20714 10792 20720 10804
rect 20027 10764 20720 10792
rect 20027 10761 20039 10764
rect 19981 10755 20039 10761
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 20898 10752 20904 10804
rect 20956 10792 20962 10804
rect 21545 10795 21603 10801
rect 21545 10792 21557 10795
rect 20956 10764 21557 10792
rect 20956 10752 20962 10764
rect 21545 10761 21557 10764
rect 21591 10792 21603 10795
rect 22554 10792 22560 10804
rect 21591 10764 22560 10792
rect 21591 10761 21603 10764
rect 21545 10755 21603 10761
rect 22554 10752 22560 10764
rect 22612 10752 22618 10804
rect 22830 10752 22836 10804
rect 22888 10752 22894 10804
rect 16485 10727 16543 10733
rect 16485 10693 16497 10727
rect 16531 10724 16543 10727
rect 21361 10727 21419 10733
rect 16531 10696 16712 10724
rect 16531 10693 16543 10696
rect 16485 10687 16543 10693
rect 14918 10656 14924 10668
rect 13924 10628 14924 10656
rect 13924 10597 13952 10628
rect 14384 10597 14412 10628
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 16684 10665 16712 10696
rect 21361 10693 21373 10727
rect 21407 10724 21419 10727
rect 21726 10724 21732 10736
rect 21407 10696 21732 10724
rect 21407 10693 21419 10696
rect 21361 10687 21419 10693
rect 21726 10684 21732 10696
rect 21784 10684 21790 10736
rect 15013 10659 15071 10665
rect 15013 10625 15025 10659
rect 15059 10656 15071 10659
rect 16669 10659 16727 10665
rect 15059 10628 16252 10656
rect 15059 10625 15071 10628
rect 15013 10619 15071 10625
rect 16224 10600 16252 10628
rect 16669 10625 16681 10659
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 18509 10659 18567 10665
rect 18509 10625 18521 10659
rect 18555 10656 18567 10659
rect 18690 10656 18696 10668
rect 18555 10628 18696 10656
rect 18555 10625 18567 10628
rect 18509 10619 18567 10625
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 12713 10591 12771 10597
rect 12400 10548 12434 10588
rect 12713 10557 12725 10591
rect 12759 10557 12771 10591
rect 12713 10551 12771 10557
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 13081 10591 13139 10597
rect 13081 10557 13093 10591
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 13265 10591 13323 10597
rect 13265 10557 13277 10591
rect 13311 10588 13323 10591
rect 13909 10591 13967 10597
rect 13909 10588 13921 10591
rect 13311 10560 13921 10588
rect 13311 10557 13323 10560
rect 13265 10551 13323 10557
rect 13909 10557 13921 10560
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 14093 10591 14151 10597
rect 14093 10557 14105 10591
rect 14139 10588 14151 10591
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 14139 10560 14289 10588
rect 14139 10557 14151 10560
rect 14093 10551 14151 10557
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 14369 10591 14427 10597
rect 14369 10557 14381 10591
rect 14415 10557 14427 10591
rect 14369 10551 14427 10557
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10588 14703 10591
rect 14826 10588 14832 10600
rect 14691 10560 14832 10588
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 12124 10492 12296 10520
rect 12406 10520 12434 10548
rect 12912 10520 12940 10551
rect 12406 10492 12940 10520
rect 14292 10520 14320 10551
rect 14660 10520 14688 10551
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 15102 10548 15108 10600
rect 15160 10548 15166 10600
rect 16206 10548 16212 10600
rect 16264 10548 16270 10600
rect 16301 10591 16359 10597
rect 16301 10557 16313 10591
rect 16347 10588 16359 10591
rect 16390 10588 16396 10600
rect 16347 10560 16396 10588
rect 16347 10557 16359 10560
rect 16301 10551 16359 10557
rect 16390 10548 16396 10560
rect 16448 10548 16454 10600
rect 16485 10591 16543 10597
rect 16485 10557 16497 10591
rect 16531 10588 16543 10591
rect 16531 10560 16804 10588
rect 16531 10557 16543 10560
rect 16485 10551 16543 10557
rect 14292 10492 14688 10520
rect 12124 10480 12130 10492
rect 16574 10480 16580 10532
rect 16632 10480 16638 10532
rect 16776 10520 16804 10560
rect 16850 10548 16856 10600
rect 16908 10548 16914 10600
rect 18230 10548 18236 10600
rect 18288 10597 18294 10600
rect 18288 10588 18300 10597
rect 18288 10560 18333 10588
rect 18288 10551 18300 10560
rect 18288 10548 18294 10551
rect 23014 10548 23020 10600
rect 23072 10548 23078 10600
rect 17770 10520 17776 10532
rect 16776 10492 17776 10520
rect 16868 10464 16896 10492
rect 17770 10480 17776 10492
rect 17828 10480 17834 10532
rect 19978 10529 19984 10532
rect 19965 10523 19984 10529
rect 19965 10489 19977 10523
rect 19965 10483 19984 10489
rect 19978 10480 19984 10483
rect 20036 10480 20042 10532
rect 20162 10480 20168 10532
rect 20220 10480 20226 10532
rect 21082 10480 21088 10532
rect 21140 10520 21146 10532
rect 21513 10523 21571 10529
rect 21513 10520 21525 10523
rect 21140 10492 21525 10520
rect 21140 10480 21146 10492
rect 21513 10489 21525 10492
rect 21559 10489 21571 10523
rect 21513 10483 21571 10489
rect 21634 10480 21640 10532
rect 21692 10520 21698 10532
rect 21729 10523 21787 10529
rect 21729 10520 21741 10523
rect 21692 10492 21741 10520
rect 21692 10480 21698 10492
rect 21729 10489 21741 10492
rect 21775 10489 21787 10523
rect 21729 10483 21787 10489
rect 8904 10424 9628 10452
rect 11977 10455 12035 10461
rect 8904 10412 8910 10424
rect 11977 10421 11989 10455
rect 12023 10452 12035 10455
rect 12434 10452 12440 10464
rect 12023 10424 12440 10452
rect 12023 10421 12035 10424
rect 11977 10415 12035 10421
rect 12434 10412 12440 10424
rect 12492 10412 12498 10464
rect 12802 10412 12808 10464
rect 12860 10412 12866 10464
rect 13265 10455 13323 10461
rect 13265 10421 13277 10455
rect 13311 10452 13323 10455
rect 13630 10452 13636 10464
rect 13311 10424 13636 10452
rect 13311 10421 13323 10424
rect 13265 10415 13323 10421
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 14001 10455 14059 10461
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 14182 10452 14188 10464
rect 14047 10424 14188 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 14553 10455 14611 10461
rect 14553 10421 14565 10455
rect 14599 10452 14611 10455
rect 14734 10452 14740 10464
rect 14599 10424 14740 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 16850 10412 16856 10464
rect 16908 10412 16914 10464
rect 17037 10455 17095 10461
rect 17037 10421 17049 10455
rect 17083 10452 17095 10455
rect 18966 10452 18972 10464
rect 17083 10424 18972 10452
rect 17083 10421 17095 10424
rect 17037 10415 17095 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 22462 10452 22468 10464
rect 22152 10424 22468 10452
rect 22152 10412 22158 10424
rect 22462 10412 22468 10424
rect 22520 10412 22526 10464
rect 552 10362 23368 10384
rect 552 10310 4322 10362
rect 4374 10310 4386 10362
rect 4438 10310 4450 10362
rect 4502 10310 4514 10362
rect 4566 10310 4578 10362
rect 4630 10310 23368 10362
rect 552 10288 23368 10310
rect 6362 10208 6368 10260
rect 6420 10208 6426 10260
rect 7282 10208 7288 10260
rect 7340 10257 7346 10260
rect 7340 10251 7359 10257
rect 7347 10248 7359 10251
rect 8846 10248 8852 10260
rect 7347 10220 7604 10248
rect 7347 10217 7359 10220
rect 7340 10211 7359 10217
rect 7340 10208 7346 10211
rect 3510 10140 3516 10192
rect 3568 10180 3574 10192
rect 3849 10183 3907 10189
rect 3849 10180 3861 10183
rect 3568 10152 3861 10180
rect 3568 10140 3574 10152
rect 3849 10149 3861 10152
rect 3895 10149 3907 10183
rect 3849 10143 3907 10149
rect 4065 10183 4123 10189
rect 4065 10149 4077 10183
rect 4111 10180 4123 10183
rect 4154 10180 4160 10192
rect 4111 10152 4160 10180
rect 4111 10149 4123 10152
rect 4065 10143 4123 10149
rect 4154 10140 4160 10152
rect 4212 10180 4218 10192
rect 4341 10183 4399 10189
rect 4341 10180 4353 10183
rect 4212 10152 4353 10180
rect 4212 10140 4218 10152
rect 4341 10149 4353 10152
rect 4387 10149 4399 10183
rect 4341 10143 4399 10149
rect 5442 10140 5448 10192
rect 5500 10180 5506 10192
rect 7101 10183 7159 10189
rect 5500 10152 6040 10180
rect 5500 10140 5506 10152
rect 4982 10072 4988 10124
rect 5040 10072 5046 10124
rect 5169 10115 5227 10121
rect 5169 10081 5181 10115
rect 5215 10081 5227 10115
rect 5169 10075 5227 10081
rect 5184 10044 5212 10075
rect 5258 10072 5264 10124
rect 5316 10072 5322 10124
rect 5350 10072 5356 10124
rect 5408 10072 5414 10124
rect 5534 10072 5540 10124
rect 5592 10072 5598 10124
rect 6012 10121 6040 10152
rect 7101 10149 7113 10183
rect 7147 10149 7159 10183
rect 7101 10143 7159 10149
rect 5997 10115 6055 10121
rect 5997 10081 6009 10115
rect 6043 10112 6055 10115
rect 6546 10112 6552 10124
rect 6043 10084 6552 10112
rect 6043 10081 6055 10084
rect 5997 10075 6055 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 5552 10044 5580 10072
rect 5184 10016 5580 10044
rect 5626 10004 5632 10056
rect 5684 10044 5690 10056
rect 5905 10047 5963 10053
rect 5905 10044 5917 10047
rect 5684 10016 5917 10044
rect 5684 10004 5690 10016
rect 5905 10013 5917 10016
rect 5951 10013 5963 10047
rect 7116 10044 7144 10143
rect 7576 10121 7604 10220
rect 8220 10220 8852 10248
rect 7561 10115 7619 10121
rect 7561 10081 7573 10115
rect 7607 10081 7619 10115
rect 7561 10075 7619 10081
rect 7650 10072 7656 10124
rect 7708 10072 7714 10124
rect 7837 10115 7895 10121
rect 7837 10081 7849 10115
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 7852 10044 7880 10075
rect 7926 10072 7932 10124
rect 7984 10112 7990 10124
rect 8220 10121 8248 10220
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 12342 10208 12348 10260
rect 12400 10208 12406 10260
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 17497 10251 17555 10257
rect 17497 10248 17509 10251
rect 17276 10220 17509 10248
rect 17276 10208 17282 10220
rect 17497 10217 17509 10220
rect 17543 10217 17555 10251
rect 17497 10211 17555 10217
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 9185 10183 9243 10189
rect 9185 10180 9197 10183
rect 8536 10152 9197 10180
rect 8536 10140 8542 10152
rect 9185 10149 9197 10152
rect 9231 10149 9243 10183
rect 9185 10143 9243 10149
rect 9398 10140 9404 10192
rect 9456 10140 9462 10192
rect 11514 10140 11520 10192
rect 11572 10180 11578 10192
rect 12360 10180 12388 10208
rect 11572 10152 12388 10180
rect 17512 10180 17540 10211
rect 17586 10208 17592 10260
rect 17644 10208 17650 10260
rect 17862 10208 17868 10260
rect 17920 10248 17926 10260
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 17920 10220 18245 10248
rect 17920 10208 17926 10220
rect 18233 10217 18245 10220
rect 18279 10217 18291 10251
rect 18233 10211 18291 10217
rect 21269 10251 21327 10257
rect 21269 10217 21281 10251
rect 21315 10248 21327 10251
rect 22094 10248 22100 10260
rect 21315 10220 22100 10248
rect 21315 10217 21327 10220
rect 21269 10211 21327 10217
rect 22094 10208 22100 10220
rect 22152 10208 22158 10260
rect 22186 10208 22192 10260
rect 22244 10248 22250 10260
rect 22373 10251 22431 10257
rect 22373 10248 22385 10251
rect 22244 10220 22385 10248
rect 22244 10208 22250 10220
rect 22373 10217 22385 10220
rect 22419 10217 22431 10251
rect 22373 10211 22431 10217
rect 18049 10183 18107 10189
rect 18049 10180 18061 10183
rect 17512 10152 18061 10180
rect 11572 10140 11578 10152
rect 8205 10115 8263 10121
rect 8205 10112 8217 10115
rect 7984 10084 8217 10112
rect 7984 10072 7990 10084
rect 8205 10081 8217 10084
rect 8251 10081 8263 10115
rect 8938 10112 8944 10124
rect 8205 10075 8263 10081
rect 8312 10084 8944 10112
rect 8110 10044 8116 10056
rect 7116 10016 8116 10044
rect 5905 10007 5963 10013
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 3697 9979 3755 9985
rect 3697 9945 3709 9979
rect 3743 9976 3755 9979
rect 4062 9976 4068 9988
rect 3743 9948 4068 9976
rect 3743 9945 3755 9948
rect 3697 9939 3755 9945
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 4709 9979 4767 9985
rect 4709 9945 4721 9979
rect 4755 9976 4767 9979
rect 6362 9976 6368 9988
rect 4755 9948 6368 9976
rect 4755 9945 4767 9948
rect 4709 9939 4767 9945
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 7650 9976 7656 9988
rect 7300 9948 7656 9976
rect 3326 9868 3332 9920
rect 3384 9908 3390 9920
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3384 9880 3893 9908
rect 3384 9868 3390 9880
rect 3881 9877 3893 9880
rect 3927 9877 3939 9911
rect 3881 9871 3939 9877
rect 4157 9911 4215 9917
rect 4157 9877 4169 9911
rect 4203 9908 4215 9911
rect 4246 9908 4252 9920
rect 4203 9880 4252 9908
rect 4203 9877 4215 9880
rect 4157 9871 4215 9877
rect 4246 9868 4252 9880
rect 4304 9868 4310 9920
rect 4341 9911 4399 9917
rect 4341 9877 4353 9911
rect 4387 9908 4399 9911
rect 4801 9911 4859 9917
rect 4801 9908 4813 9911
rect 4387 9880 4813 9908
rect 4387 9877 4399 9880
rect 4341 9871 4399 9877
rect 4801 9877 4813 9880
rect 4847 9877 4859 9911
rect 4801 9871 4859 9877
rect 5445 9911 5503 9917
rect 5445 9877 5457 9911
rect 5491 9908 5503 9911
rect 5994 9908 6000 9920
rect 5491 9880 6000 9908
rect 5491 9877 5503 9880
rect 5445 9871 5503 9877
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7300 9917 7328 9948
rect 7650 9936 7656 9948
rect 7708 9976 7714 9988
rect 8312 9985 8340 10084
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 11422 10072 11428 10124
rect 11480 10072 11486 10124
rect 11992 10121 12020 10152
rect 18049 10149 18061 10152
rect 18095 10149 18107 10183
rect 18049 10143 18107 10149
rect 21082 10140 21088 10192
rect 21140 10180 21146 10192
rect 22002 10180 22008 10192
rect 21140 10152 22008 10180
rect 21140 10140 21146 10152
rect 22002 10140 22008 10152
rect 22060 10180 22066 10192
rect 22281 10183 22339 10189
rect 22281 10180 22293 10183
rect 22060 10152 22293 10180
rect 22060 10140 22066 10152
rect 22281 10149 22293 10152
rect 22327 10149 22339 10183
rect 22281 10143 22339 10149
rect 11977 10115 12035 10121
rect 11977 10081 11989 10115
rect 12023 10081 12035 10115
rect 11977 10075 12035 10081
rect 12066 10072 12072 10124
rect 12124 10072 12130 10124
rect 12253 10115 12311 10121
rect 12253 10081 12265 10115
rect 12299 10112 12311 10115
rect 12345 10115 12403 10121
rect 12345 10112 12357 10115
rect 12299 10084 12357 10112
rect 12299 10081 12311 10084
rect 12253 10075 12311 10081
rect 12345 10081 12357 10084
rect 12391 10081 12403 10115
rect 12345 10075 12403 10081
rect 12529 10115 12587 10121
rect 12529 10081 12541 10115
rect 12575 10112 12587 10115
rect 12802 10112 12808 10124
rect 12575 10084 12808 10112
rect 12575 10081 12587 10084
rect 12529 10075 12587 10081
rect 8481 10047 8539 10053
rect 8481 10013 8493 10047
rect 8527 10044 8539 10047
rect 8570 10044 8576 10056
rect 8527 10016 8576 10044
rect 8527 10013 8539 10016
rect 8481 10007 8539 10013
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 8846 10004 8852 10056
rect 8904 10004 8910 10056
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 8297 9979 8355 9985
rect 8297 9976 8309 9979
rect 7708 9948 8309 9976
rect 7708 9936 7714 9948
rect 8297 9945 8309 9948
rect 8343 9945 8355 9979
rect 11532 9976 11560 10007
rect 12544 9976 12572 10075
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 14274 10072 14280 10124
rect 14332 10072 14338 10124
rect 14734 10072 14740 10124
rect 14792 10072 14798 10124
rect 14921 10115 14979 10121
rect 14921 10081 14933 10115
rect 14967 10081 14979 10115
rect 14921 10075 14979 10081
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 14936 10044 14964 10075
rect 16942 10072 16948 10124
rect 17000 10112 17006 10124
rect 17221 10115 17279 10121
rect 17221 10112 17233 10115
rect 17000 10084 17233 10112
rect 17000 10072 17006 10084
rect 17221 10081 17233 10084
rect 17267 10081 17279 10115
rect 17221 10075 17279 10081
rect 17402 10072 17408 10124
rect 17460 10072 17466 10124
rect 17770 10072 17776 10124
rect 17828 10072 17834 10124
rect 17862 10072 17868 10124
rect 17920 10072 17926 10124
rect 20714 10072 20720 10124
rect 20772 10072 20778 10124
rect 20898 10072 20904 10124
rect 20956 10072 20962 10124
rect 21174 10072 21180 10124
rect 21232 10112 21238 10124
rect 21634 10112 21640 10124
rect 21232 10084 21640 10112
rect 21232 10072 21238 10084
rect 21634 10072 21640 10084
rect 21692 10112 21698 10124
rect 22097 10115 22155 10121
rect 22097 10112 22109 10115
rect 21692 10084 22109 10112
rect 21692 10072 21698 10084
rect 22097 10081 22109 10084
rect 22143 10081 22155 10115
rect 22097 10075 22155 10081
rect 14240 10016 14964 10044
rect 14240 10004 14246 10016
rect 21450 10004 21456 10056
rect 21508 10004 21514 10056
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10013 21603 10047
rect 21545 10007 21603 10013
rect 21729 10047 21787 10053
rect 21729 10013 21741 10047
rect 21775 10013 21787 10047
rect 22112 10044 22140 10075
rect 22738 10072 22744 10124
rect 22796 10072 22802 10124
rect 22649 10047 22707 10053
rect 22649 10044 22661 10047
rect 22112 10016 22661 10044
rect 21729 10007 21787 10013
rect 22649 10013 22661 10016
rect 22695 10044 22707 10047
rect 22830 10044 22836 10056
rect 22695 10016 22836 10044
rect 22695 10013 22707 10016
rect 22649 10007 22707 10013
rect 8297 9939 8355 9945
rect 8588 9948 9260 9976
rect 11532 9948 12572 9976
rect 14645 9979 14703 9985
rect 8588 9920 8616 9948
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 7064 9880 7297 9908
rect 7064 9868 7070 9880
rect 7285 9877 7297 9880
rect 7331 9877 7343 9911
rect 7285 9871 7343 9877
rect 7466 9868 7472 9920
rect 7524 9868 7530 9920
rect 7834 9868 7840 9920
rect 7892 9868 7898 9920
rect 8570 9868 8576 9920
rect 8628 9868 8634 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8720 9880 8769 9908
rect 8720 9868 8726 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 9033 9911 9091 9917
rect 9033 9877 9045 9911
rect 9079 9908 9091 9911
rect 9122 9908 9128 9920
rect 9079 9880 9128 9908
rect 9079 9877 9091 9880
rect 9033 9871 9091 9877
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 9232 9917 9260 9948
rect 14645 9945 14657 9979
rect 14691 9976 14703 9979
rect 14918 9976 14924 9988
rect 14691 9948 14924 9976
rect 14691 9945 14703 9948
rect 14645 9939 14703 9945
rect 14918 9936 14924 9948
rect 14976 9936 14982 9988
rect 16666 9936 16672 9988
rect 16724 9976 16730 9988
rect 17586 9976 17592 9988
rect 16724 9948 17592 9976
rect 16724 9936 16730 9948
rect 17586 9936 17592 9948
rect 17644 9936 17650 9988
rect 20806 9936 20812 9988
rect 20864 9976 20870 9988
rect 21560 9976 21588 10007
rect 20864 9948 21588 9976
rect 21744 9976 21772 10007
rect 22830 10004 22836 10016
rect 22888 10004 22894 10056
rect 21744 9948 22094 9976
rect 20864 9936 20870 9948
rect 9217 9911 9275 9917
rect 9217 9877 9229 9911
rect 9263 9908 9275 9911
rect 9306 9908 9312 9920
rect 9263 9880 9312 9908
rect 9263 9877 9275 9880
rect 9217 9871 9275 9877
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 11698 9868 11704 9920
rect 11756 9868 11762 9920
rect 12342 9868 12348 9920
rect 12400 9868 12406 9920
rect 14458 9868 14464 9920
rect 14516 9908 14522 9920
rect 14737 9911 14795 9917
rect 14737 9908 14749 9911
rect 14516 9880 14749 9908
rect 14516 9868 14522 9880
rect 14737 9877 14749 9880
rect 14783 9877 14795 9911
rect 14737 9871 14795 9877
rect 21085 9911 21143 9917
rect 21085 9877 21097 9911
rect 21131 9908 21143 9911
rect 21266 9908 21272 9920
rect 21131 9880 21272 9908
rect 21131 9877 21143 9880
rect 21085 9871 21143 9877
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 21358 9868 21364 9920
rect 21416 9908 21422 9920
rect 21913 9911 21971 9917
rect 21913 9908 21925 9911
rect 21416 9880 21925 9908
rect 21416 9868 21422 9880
rect 21913 9877 21925 9880
rect 21959 9877 21971 9911
rect 22066 9908 22094 9948
rect 22370 9908 22376 9920
rect 22066 9880 22376 9908
rect 21913 9871 21971 9877
rect 22370 9868 22376 9880
rect 22428 9868 22434 9920
rect 22554 9868 22560 9920
rect 22612 9868 22618 9920
rect 552 9818 23368 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 23368 9818
rect 552 9744 23368 9766
rect 3326 9664 3332 9716
rect 3384 9664 3390 9716
rect 3510 9664 3516 9716
rect 3568 9704 3574 9716
rect 3881 9707 3939 9713
rect 3881 9704 3893 9707
rect 3568 9676 3893 9704
rect 3568 9664 3574 9676
rect 3881 9673 3893 9676
rect 3927 9673 3939 9707
rect 3881 9667 3939 9673
rect 4982 9664 4988 9716
rect 5040 9704 5046 9716
rect 5353 9707 5411 9713
rect 5353 9704 5365 9707
rect 5040 9676 5365 9704
rect 5040 9664 5046 9676
rect 5353 9673 5365 9676
rect 5399 9704 5411 9707
rect 5442 9704 5448 9716
rect 5399 9676 5448 9704
rect 5399 9673 5411 9676
rect 5353 9667 5411 9673
rect 5442 9664 5448 9676
rect 5500 9664 5506 9716
rect 5813 9707 5871 9713
rect 5813 9673 5825 9707
rect 5859 9704 5871 9707
rect 6089 9707 6147 9713
rect 6089 9704 6101 9707
rect 5859 9676 6101 9704
rect 5859 9673 5871 9676
rect 5813 9667 5871 9673
rect 6089 9673 6101 9676
rect 6135 9673 6147 9707
rect 6089 9667 6147 9673
rect 6546 9664 6552 9716
rect 6604 9664 6610 9716
rect 7469 9707 7527 9713
rect 7469 9673 7481 9707
rect 7515 9704 7527 9707
rect 7834 9704 7840 9716
rect 7515 9676 7840 9704
rect 7515 9673 7527 9676
rect 7469 9667 7527 9673
rect 7834 9664 7840 9676
rect 7892 9664 7898 9716
rect 8846 9664 8852 9716
rect 8904 9664 8910 9716
rect 14645 9707 14703 9713
rect 14645 9673 14657 9707
rect 14691 9704 14703 9707
rect 15473 9707 15531 9713
rect 15473 9704 15485 9707
rect 14691 9676 15485 9704
rect 14691 9673 14703 9676
rect 14645 9667 14703 9673
rect 15473 9673 15485 9676
rect 15519 9673 15531 9707
rect 15473 9667 15531 9673
rect 16666 9664 16672 9716
rect 16724 9664 16730 9716
rect 18969 9707 19027 9713
rect 18969 9673 18981 9707
rect 19015 9704 19027 9707
rect 19245 9707 19303 9713
rect 19245 9704 19257 9707
rect 19015 9676 19257 9704
rect 19015 9673 19027 9676
rect 18969 9667 19027 9673
rect 19245 9673 19257 9676
rect 19291 9673 19303 9707
rect 19245 9667 19303 9673
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 21177 9707 21235 9713
rect 20772 9676 20852 9704
rect 20772 9664 20778 9676
rect 5905 9639 5963 9645
rect 5905 9605 5917 9639
rect 5951 9605 5963 9639
rect 5905 9599 5963 9605
rect 5920 9568 5948 9599
rect 6362 9596 6368 9648
rect 6420 9596 6426 9648
rect 8202 9596 8208 9648
rect 8260 9596 8266 9648
rect 8864 9636 8892 9664
rect 8772 9608 8892 9636
rect 14093 9639 14151 9645
rect 6086 9568 6092 9580
rect 5920 9540 6092 9568
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 8352 9540 8401 9568
rect 8352 9528 8358 9540
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 3237 9503 3295 9509
rect 3237 9469 3249 9503
rect 3283 9469 3295 9503
rect 3237 9463 3295 9469
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9500 3479 9503
rect 3467 9472 3740 9500
rect 3467 9469 3479 9472
rect 3421 9463 3479 9469
rect 3252 9432 3280 9463
rect 3712 9441 3740 9472
rect 3970 9460 3976 9512
rect 4028 9460 4034 9512
rect 4246 9509 4252 9512
rect 4240 9500 4252 9509
rect 4207 9472 4252 9500
rect 4240 9463 4252 9472
rect 4246 9460 4252 9463
rect 4304 9460 4310 9512
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 5408 9472 5457 9500
rect 5408 9460 5414 9472
rect 5445 9469 5457 9472
rect 5491 9469 5503 9503
rect 5445 9463 5503 9469
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 5592 9472 5641 9500
rect 5592 9460 5598 9472
rect 5629 9469 5641 9472
rect 5675 9500 5687 9503
rect 5675 9472 6776 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 3513 9435 3571 9441
rect 3513 9432 3525 9435
rect 3252 9404 3525 9432
rect 3513 9401 3525 9404
rect 3559 9401 3571 9435
rect 3513 9395 3571 9401
rect 3697 9435 3755 9441
rect 3697 9401 3709 9435
rect 3743 9432 3755 9435
rect 5552 9432 5580 9460
rect 3743 9404 5580 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 3528 9364 3556 9395
rect 5994 9392 6000 9444
rect 6052 9441 6058 9444
rect 6748 9441 6776 9472
rect 7190 9460 7196 9512
rect 7248 9500 7254 9512
rect 7285 9503 7343 9509
rect 7285 9500 7297 9503
rect 7248 9472 7297 9500
rect 7248 9460 7254 9472
rect 7285 9469 7297 9472
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 7466 9460 7472 9512
rect 7524 9460 7530 9512
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9469 7987 9503
rect 7929 9463 7987 9469
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8570 9500 8576 9512
rect 8067 9472 8576 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 6052 9435 6115 9441
rect 6052 9401 6069 9435
rect 6103 9401 6115 9435
rect 6052 9395 6115 9401
rect 6273 9435 6331 9441
rect 6273 9401 6285 9435
rect 6319 9432 6331 9435
rect 6517 9435 6575 9441
rect 6517 9432 6529 9435
rect 6319 9404 6529 9432
rect 6319 9401 6331 9404
rect 6273 9395 6331 9401
rect 6517 9401 6529 9404
rect 6563 9401 6575 9435
rect 6517 9395 6575 9401
rect 6733 9435 6791 9441
rect 6733 9401 6745 9435
rect 6779 9401 6791 9435
rect 6733 9395 6791 9401
rect 6052 9392 6058 9395
rect 5258 9364 5264 9376
rect 3528 9336 5264 9364
rect 5258 9324 5264 9336
rect 5316 9364 5322 9376
rect 5442 9364 5448 9376
rect 5316 9336 5448 9364
rect 5316 9324 5322 9336
rect 5442 9324 5448 9336
rect 5500 9364 5506 9376
rect 6288 9364 6316 9395
rect 5500 9336 6316 9364
rect 5500 9324 5506 9336
rect 7650 9324 7656 9376
rect 7708 9324 7714 9376
rect 7944 9364 7972 9463
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8772 9509 8800 9608
rect 14093 9605 14105 9639
rect 14139 9636 14151 9639
rect 15933 9639 15991 9645
rect 14139 9608 15608 9636
rect 14139 9605 14151 9608
rect 14093 9599 14151 9605
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9568 8907 9571
rect 8938 9568 8944 9580
rect 8895 9540 8944 9568
rect 8895 9537 8907 9540
rect 8849 9531 8907 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 9306 9528 9312 9580
rect 9364 9528 9370 9580
rect 11425 9571 11483 9577
rect 11425 9537 11437 9571
rect 11471 9568 11483 9571
rect 12342 9568 12348 9580
rect 11471 9540 12348 9568
rect 11471 9537 11483 9540
rect 11425 9531 11483 9537
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 13630 9528 13636 9580
rect 13688 9528 13694 9580
rect 14458 9528 14464 9580
rect 14516 9528 14522 9580
rect 14918 9528 14924 9580
rect 14976 9528 14982 9580
rect 15580 9577 15608 9608
rect 15933 9605 15945 9639
rect 15979 9636 15991 9639
rect 16574 9636 16580 9648
rect 15979 9608 16580 9636
rect 15979 9605 15991 9608
rect 15933 9599 15991 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 20824 9645 20852 9676
rect 21177 9673 21189 9707
rect 21223 9704 21235 9707
rect 21358 9704 21364 9716
rect 21223 9676 21364 9704
rect 21223 9673 21235 9676
rect 21177 9667 21235 9673
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 22830 9664 22836 9716
rect 22888 9664 22894 9716
rect 20809 9639 20867 9645
rect 20809 9605 20821 9639
rect 20855 9605 20867 9639
rect 20809 9599 20867 9605
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 16132 9540 16804 9568
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9469 8815 9503
rect 8757 9463 8815 9469
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 9490 9500 9496 9512
rect 9447 9472 9496 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 11330 9460 11336 9512
rect 11388 9460 11394 9512
rect 13722 9460 13728 9512
rect 13780 9460 13786 9512
rect 14366 9460 14372 9512
rect 14424 9460 14430 9512
rect 15013 9503 15071 9509
rect 15013 9469 15025 9503
rect 15059 9500 15071 9503
rect 15194 9500 15200 9512
rect 15059 9472 15200 9500
rect 15059 9469 15071 9472
rect 15013 9463 15071 9469
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 16132 9509 16160 9540
rect 15749 9503 15807 9509
rect 15749 9500 15761 9503
rect 15396 9472 15761 9500
rect 8205 9435 8263 9441
rect 8205 9401 8217 9435
rect 8251 9432 8263 9435
rect 8251 9404 8616 9432
rect 8251 9401 8263 9404
rect 8205 9395 8263 9401
rect 8588 9376 8616 9404
rect 8478 9364 8484 9376
rect 7944 9336 8484 9364
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 8570 9324 8576 9376
rect 8628 9364 8634 9376
rect 9398 9364 9404 9376
rect 8628 9336 9404 9364
rect 8628 9324 8634 9336
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 11054 9364 11060 9376
rect 9815 9336 11060 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 11701 9367 11759 9373
rect 11701 9333 11713 9367
rect 11747 9364 11759 9367
rect 12250 9364 12256 9376
rect 11747 9336 12256 9364
rect 11747 9333 11759 9336
rect 11701 9327 11759 9333
rect 12250 9324 12256 9336
rect 12308 9324 12314 9376
rect 15396 9373 15424 9472
rect 15749 9469 15761 9472
rect 15795 9469 15807 9503
rect 15749 9463 15807 9469
rect 16117 9503 16175 9509
rect 16117 9469 16129 9503
rect 16163 9469 16175 9503
rect 16117 9463 16175 9469
rect 16393 9503 16451 9509
rect 16393 9469 16405 9503
rect 16439 9500 16451 9503
rect 16666 9500 16672 9512
rect 16439 9472 16672 9500
rect 16439 9469 16451 9472
rect 16393 9463 16451 9469
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 16776 9500 16804 9540
rect 18046 9528 18052 9580
rect 18104 9568 18110 9580
rect 18690 9568 18696 9580
rect 18104 9540 18696 9568
rect 18104 9528 18110 9540
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 20349 9571 20407 9577
rect 20349 9537 20361 9571
rect 20395 9568 20407 9571
rect 21174 9568 21180 9580
rect 20395 9540 21180 9568
rect 20395 9537 20407 9540
rect 20349 9531 20407 9537
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 17402 9500 17408 9512
rect 16776 9472 17408 9500
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9500 19487 9503
rect 20533 9503 20591 9509
rect 19475 9472 19739 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 15470 9392 15476 9444
rect 15528 9392 15534 9444
rect 16209 9435 16267 9441
rect 16209 9401 16221 9435
rect 16255 9432 16267 9435
rect 16255 9404 16712 9432
rect 16255 9401 16267 9404
rect 16209 9395 16267 9401
rect 15381 9367 15439 9373
rect 15381 9333 15393 9367
rect 15427 9333 15439 9367
rect 15381 9327 15439 9333
rect 16574 9324 16580 9376
rect 16632 9324 16638 9376
rect 16684 9364 16712 9404
rect 16758 9392 16764 9444
rect 16816 9432 16822 9444
rect 17782 9435 17840 9441
rect 17782 9432 17794 9435
rect 16816 9404 17794 9432
rect 16816 9392 16822 9404
rect 17782 9401 17794 9404
rect 17828 9401 17840 9435
rect 17782 9395 17840 9401
rect 19150 9392 19156 9444
rect 19208 9392 19214 9444
rect 19610 9392 19616 9444
rect 19668 9392 19674 9444
rect 19711 9432 19739 9472
rect 20533 9469 20545 9503
rect 20579 9500 20591 9503
rect 21082 9500 21088 9512
rect 20579 9472 21088 9500
rect 20579 9469 20591 9472
rect 20533 9463 20591 9469
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 21358 9460 21364 9512
rect 21416 9500 21422 9512
rect 21453 9503 21511 9509
rect 21453 9500 21465 9503
rect 21416 9472 21465 9500
rect 21416 9460 21422 9472
rect 21453 9469 21465 9472
rect 21499 9500 21511 9503
rect 21542 9500 21548 9512
rect 21499 9472 21548 9500
rect 21499 9469 21511 9472
rect 21453 9463 21511 9469
rect 21542 9460 21548 9472
rect 21600 9500 21606 9512
rect 21600 9472 21864 9500
rect 21600 9460 21606 9472
rect 21836 9444 21864 9472
rect 19886 9432 19892 9444
rect 19711 9404 19892 9432
rect 19886 9392 19892 9404
rect 19944 9432 19950 9444
rect 20806 9432 20812 9444
rect 19944 9404 20812 9432
rect 19944 9392 19950 9404
rect 20806 9392 20812 9404
rect 20864 9392 20870 9444
rect 21698 9435 21756 9441
rect 21698 9432 21710 9435
rect 21376 9404 21710 9432
rect 16850 9364 16856 9376
rect 16684 9336 16856 9364
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 18782 9324 18788 9376
rect 18840 9324 18846 9376
rect 18953 9367 19011 9373
rect 18953 9333 18965 9367
rect 18999 9364 19011 9367
rect 19518 9364 19524 9376
rect 18999 9336 19524 9364
rect 18999 9333 19011 9336
rect 18953 9327 19011 9333
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 21376 9373 21404 9404
rect 21698 9401 21710 9404
rect 21744 9401 21756 9435
rect 21698 9395 21756 9401
rect 21818 9392 21824 9444
rect 21876 9392 21882 9444
rect 21177 9367 21235 9373
rect 21177 9364 21189 9367
rect 21140 9336 21189 9364
rect 21140 9324 21146 9336
rect 21177 9333 21189 9336
rect 21223 9333 21235 9367
rect 21177 9327 21235 9333
rect 21361 9367 21419 9373
rect 21361 9333 21373 9367
rect 21407 9333 21419 9367
rect 21361 9327 21419 9333
rect 552 9274 23368 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 23368 9274
rect 552 9200 23368 9222
rect 4982 9120 4988 9172
rect 5040 9160 5046 9172
rect 5261 9163 5319 9169
rect 5261 9160 5273 9163
rect 5040 9132 5273 9160
rect 5040 9120 5046 9132
rect 5261 9129 5273 9132
rect 5307 9129 5319 9163
rect 5261 9123 5319 9129
rect 7193 9163 7251 9169
rect 7193 9129 7205 9163
rect 7239 9129 7251 9163
rect 7193 9123 7251 9129
rect 9401 9163 9459 9169
rect 9401 9129 9413 9163
rect 9447 9160 9459 9163
rect 12713 9163 12771 9169
rect 9447 9132 12296 9160
rect 9447 9129 9459 9132
rect 9401 9123 9459 9129
rect 3872 9095 3930 9101
rect 3872 9061 3884 9095
rect 3918 9092 3930 9095
rect 4062 9092 4068 9104
rect 3918 9064 4068 9092
rect 3918 9061 3930 9064
rect 3872 9055 3930 9061
rect 4062 9052 4068 9064
rect 4120 9052 4126 9104
rect 5074 9052 5080 9104
rect 5132 9092 5138 9104
rect 5353 9095 5411 9101
rect 5353 9092 5365 9095
rect 5132 9064 5365 9092
rect 5132 9052 5138 9064
rect 5353 9061 5365 9064
rect 5399 9092 5411 9095
rect 7098 9092 7104 9104
rect 5399 9064 7104 9092
rect 5399 9061 5411 9064
rect 5353 9055 5411 9061
rect 7098 9052 7104 9064
rect 7156 9092 7162 9104
rect 7208 9092 7236 9123
rect 7156 9064 7236 9092
rect 7156 9052 7162 9064
rect 7650 9052 7656 9104
rect 7708 9092 7714 9104
rect 12268 9101 12296 9132
rect 12713 9129 12725 9163
rect 12759 9160 12771 9163
rect 15470 9160 15476 9172
rect 12759 9132 15476 9160
rect 12759 9129 12771 9132
rect 12713 9123 12771 9129
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 16758 9120 16764 9172
rect 16816 9120 16822 9172
rect 17310 9120 17316 9172
rect 17368 9120 17374 9172
rect 19886 9120 19892 9172
rect 19944 9160 19950 9172
rect 19944 9132 20024 9160
rect 19944 9120 19950 9132
rect 8941 9095 8999 9101
rect 8941 9092 8953 9095
rect 7708 9064 8953 9092
rect 7708 9052 7714 9064
rect 8941 9061 8953 9064
rect 8987 9061 8999 9095
rect 8941 9055 8999 9061
rect 12253 9095 12311 9101
rect 12253 9061 12265 9095
rect 12299 9061 12311 9095
rect 12253 9055 12311 9061
rect 14737 9095 14795 9101
rect 14737 9061 14749 9095
rect 14783 9092 14795 9095
rect 15194 9092 15200 9104
rect 14783 9064 15200 9092
rect 14783 9061 14795 9064
rect 14737 9055 14795 9061
rect 15194 9052 15200 9064
rect 15252 9052 15258 9104
rect 16482 9052 16488 9104
rect 16540 9052 16546 9104
rect 16666 9052 16672 9104
rect 16724 9092 16730 9104
rect 16945 9095 17003 9101
rect 16945 9092 16957 9095
rect 16724 9064 16957 9092
rect 16724 9052 16730 9064
rect 16945 9061 16957 9064
rect 16991 9092 17003 9095
rect 17328 9092 17356 9120
rect 16991 9064 17356 9092
rect 16991 9061 17003 9064
rect 16945 9055 17003 9061
rect 17402 9052 17408 9104
rect 17460 9092 17466 9104
rect 17557 9095 17615 9101
rect 17557 9092 17569 9095
rect 17460 9064 17569 9092
rect 17460 9052 17466 9064
rect 17557 9061 17569 9064
rect 17603 9061 17615 9095
rect 17557 9055 17615 9061
rect 17770 9052 17776 9104
rect 17828 9052 17834 9104
rect 18782 9101 18788 9104
rect 18776 9092 18788 9101
rect 18743 9064 18788 9092
rect 18776 9055 18788 9064
rect 18782 9052 18788 9055
rect 18840 9052 18846 9104
rect 19426 9052 19432 9104
rect 19484 9052 19490 9104
rect 19996 9101 20024 9132
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 20441 9163 20499 9169
rect 20441 9160 20453 9163
rect 20404 9132 20453 9160
rect 20404 9120 20410 9132
rect 20441 9129 20453 9132
rect 20487 9129 20499 9163
rect 20898 9160 20904 9172
rect 20441 9123 20499 9129
rect 20548 9132 20904 9160
rect 20548 9101 20576 9132
rect 20898 9120 20904 9132
rect 20956 9120 20962 9172
rect 21085 9163 21143 9169
rect 21085 9129 21097 9163
rect 21131 9160 21143 9163
rect 21450 9160 21456 9172
rect 21131 9132 21456 9160
rect 21131 9129 21143 9132
rect 21085 9123 21143 9129
rect 21450 9120 21456 9132
rect 21508 9120 21514 9172
rect 22554 9120 22560 9172
rect 22612 9160 22618 9172
rect 22649 9163 22707 9169
rect 22649 9160 22661 9163
rect 22612 9132 22661 9160
rect 22612 9120 22618 9132
rect 22649 9129 22661 9132
rect 22695 9129 22707 9163
rect 22649 9123 22707 9129
rect 19981 9095 20039 9101
rect 19981 9061 19993 9095
rect 20027 9061 20039 9095
rect 19981 9055 20039 9061
rect 20533 9095 20591 9101
rect 20533 9061 20545 9095
rect 20579 9061 20591 9095
rect 20990 9092 20996 9104
rect 20533 9055 20591 9061
rect 20732 9064 20996 9092
rect 5442 8984 5448 9036
rect 5500 8984 5506 9036
rect 6086 9033 6092 9036
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 8993 5871 9027
rect 5813 8987 5871 8993
rect 6080 8987 6092 9033
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8925 3663 8959
rect 3605 8919 3663 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5534 8956 5540 8968
rect 5123 8928 5540 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 3620 8820 3648 8919
rect 4985 8891 5043 8897
rect 4985 8857 4997 8891
rect 5031 8888 5043 8891
rect 5092 8888 5120 8919
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5828 8888 5856 8987
rect 6086 8984 6092 8987
rect 6144 8984 6150 9036
rect 7926 8984 7932 9036
rect 7984 9024 7990 9036
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 7984 8996 8401 9024
rect 7984 8984 7990 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 9122 8984 9128 9036
rect 9180 9024 9186 9036
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 9180 8996 9229 9024
rect 9180 8984 9186 8996
rect 9217 8993 9229 8996
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 11146 8984 11152 9036
rect 11204 8984 11210 9036
rect 11790 8984 11796 9036
rect 11848 8984 11854 9036
rect 12529 9027 12587 9033
rect 12529 8993 12541 9027
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 8294 8916 8300 8968
rect 8352 8916 8358 8968
rect 9033 8959 9091 8965
rect 9033 8956 9045 8959
rect 8772 8928 9045 8956
rect 8772 8897 8800 8928
rect 9033 8925 9045 8928
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 11054 8916 11060 8968
rect 11112 8916 11118 8968
rect 11698 8916 11704 8968
rect 11756 8916 11762 8968
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 11900 8928 12357 8956
rect 5031 8860 5120 8888
rect 5184 8860 5856 8888
rect 5031 8857 5043 8860
rect 4985 8851 5043 8857
rect 3970 8820 3976 8832
rect 3620 8792 3976 8820
rect 3970 8780 3976 8792
rect 4028 8820 4034 8832
rect 5184 8820 5212 8860
rect 4028 8792 5212 8820
rect 4028 8780 4034 8792
rect 5626 8780 5632 8832
rect 5684 8780 5690 8832
rect 5828 8820 5856 8860
rect 8757 8891 8815 8897
rect 8757 8857 8769 8891
rect 8803 8857 8815 8891
rect 8757 8851 8815 8857
rect 11517 8891 11575 8897
rect 11517 8857 11529 8891
rect 11563 8888 11575 8891
rect 11900 8888 11928 8928
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 11563 8860 11928 8888
rect 12161 8891 12219 8897
rect 11563 8857 11575 8860
rect 11517 8851 11575 8857
rect 12161 8857 12173 8891
rect 12207 8888 12219 8891
rect 12544 8888 12572 8987
rect 14366 8984 14372 9036
rect 14424 9024 14430 9036
rect 14645 9027 14703 9033
rect 14645 9024 14657 9027
rect 14424 8996 14657 9024
rect 14424 8984 14430 8996
rect 14645 8993 14657 8996
rect 14691 8993 14703 9027
rect 14645 8987 14703 8993
rect 14829 9027 14887 9033
rect 14829 8993 14841 9027
rect 14875 8993 14887 9027
rect 14829 8987 14887 8993
rect 18509 9027 18567 9033
rect 18509 8993 18521 9027
rect 18555 9024 18567 9027
rect 18598 9024 18604 9036
rect 18555 8996 18604 9024
rect 18555 8993 18567 8996
rect 18509 8987 18567 8993
rect 14550 8916 14556 8968
rect 14608 8956 14614 8968
rect 14844 8956 14872 8987
rect 18598 8984 18604 8996
rect 18656 9024 18662 9036
rect 19444 9024 19472 9052
rect 19702 9024 19708 9036
rect 18656 8996 19708 9024
rect 18656 8984 18662 8996
rect 19702 8984 19708 8996
rect 19760 9024 19766 9036
rect 20732 9033 20760 9064
rect 20990 9052 20996 9064
rect 21048 9052 21054 9104
rect 20257 9027 20315 9033
rect 19760 8996 20024 9024
rect 19760 8984 19766 8996
rect 14608 8928 14872 8956
rect 14608 8916 14614 8928
rect 15010 8916 15016 8968
rect 15068 8956 15074 8968
rect 16298 8956 16304 8968
rect 15068 8928 16304 8956
rect 15068 8916 15074 8928
rect 16298 8916 16304 8928
rect 16356 8956 16362 8968
rect 18046 8956 18052 8968
rect 16356 8928 18052 8956
rect 16356 8916 16362 8928
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 12207 8860 12572 8888
rect 12207 8857 12219 8860
rect 12161 8851 12219 8857
rect 14458 8848 14464 8900
rect 14516 8848 14522 8900
rect 16574 8848 16580 8900
rect 16632 8888 16638 8900
rect 17313 8891 17371 8897
rect 16632 8860 16988 8888
rect 16632 8848 16638 8860
rect 6822 8820 6828 8832
rect 5828 8792 6828 8820
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8260 8792 8953 8820
rect 8260 8780 8266 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 12250 8780 12256 8832
rect 12308 8780 12314 8832
rect 15013 8823 15071 8829
rect 15013 8789 15025 8823
rect 15059 8820 15071 8823
rect 16482 8820 16488 8832
rect 15059 8792 16488 8820
rect 15059 8789 15071 8792
rect 15013 8783 15071 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 16960 8829 16988 8860
rect 17313 8857 17325 8891
rect 17359 8888 17371 8891
rect 17405 8891 17463 8897
rect 17405 8888 17417 8891
rect 17359 8860 17417 8888
rect 17359 8857 17371 8860
rect 17313 8851 17371 8857
rect 17405 8857 17417 8860
rect 17451 8888 17463 8891
rect 17862 8888 17868 8900
rect 17451 8860 17868 8888
rect 17451 8857 17463 8860
rect 17405 8851 17463 8857
rect 17862 8848 17868 8860
rect 17920 8848 17926 8900
rect 19996 8888 20024 8996
rect 20257 8993 20269 9027
rect 20303 9024 20315 9027
rect 20717 9027 20775 9033
rect 20717 9024 20729 9027
rect 20303 8996 20729 9024
rect 20303 8993 20315 8996
rect 20257 8987 20315 8993
rect 20717 8993 20729 8996
rect 20763 8993 20775 9027
rect 20717 8987 20775 8993
rect 20806 8984 20812 9036
rect 20864 8984 20870 9036
rect 20901 9027 20959 9033
rect 20901 8993 20913 9027
rect 20947 8993 20959 9027
rect 20901 8987 20959 8993
rect 20070 8916 20076 8968
rect 20128 8956 20134 8968
rect 20165 8959 20223 8965
rect 20165 8956 20177 8959
rect 20128 8928 20177 8956
rect 20128 8916 20134 8928
rect 20165 8925 20177 8928
rect 20211 8956 20223 8959
rect 20916 8956 20944 8987
rect 21174 8984 21180 9036
rect 21232 9024 21238 9036
rect 21525 9027 21583 9033
rect 21525 9024 21537 9027
rect 21232 8996 21537 9024
rect 21232 8984 21238 8996
rect 21525 8993 21537 8996
rect 21571 8993 21583 9027
rect 21525 8987 21583 8993
rect 20211 8928 20944 8956
rect 21269 8959 21327 8965
rect 20211 8925 20223 8928
rect 20165 8919 20223 8925
rect 21269 8925 21281 8959
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 21284 8888 21312 8919
rect 19996 8860 21312 8888
rect 16945 8823 17003 8829
rect 16945 8789 16957 8823
rect 16991 8789 17003 8823
rect 16945 8783 17003 8789
rect 17586 8780 17592 8832
rect 17644 8780 17650 8832
rect 20257 8823 20315 8829
rect 20257 8789 20269 8823
rect 20303 8820 20315 8823
rect 20806 8820 20812 8832
rect 20303 8792 20812 8820
rect 20303 8789 20315 8792
rect 20257 8783 20315 8789
rect 20806 8780 20812 8792
rect 20864 8780 20870 8832
rect 21284 8820 21312 8860
rect 22002 8820 22008 8832
rect 21284 8792 22008 8820
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 552 8730 23368 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 23368 8730
rect 552 8656 23368 8678
rect 5905 8619 5963 8625
rect 5905 8585 5917 8619
rect 5951 8585 5963 8619
rect 5905 8579 5963 8585
rect 5537 8551 5595 8557
rect 5537 8517 5549 8551
rect 5583 8548 5595 8551
rect 5626 8548 5632 8560
rect 5583 8520 5632 8548
rect 5583 8517 5595 8520
rect 5537 8511 5595 8517
rect 5626 8508 5632 8520
rect 5684 8508 5690 8560
rect 5920 8548 5948 8579
rect 6086 8576 6092 8628
rect 6144 8576 6150 8628
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 11057 8619 11115 8625
rect 11057 8616 11069 8619
rect 10560 8588 11069 8616
rect 10560 8576 10566 8588
rect 11057 8585 11069 8588
rect 11103 8616 11115 8619
rect 11330 8616 11336 8628
rect 11103 8588 11336 8616
rect 11103 8585 11115 8588
rect 11057 8579 11115 8585
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 13906 8576 13912 8628
rect 13964 8576 13970 8628
rect 14366 8576 14372 8628
rect 14424 8616 14430 8628
rect 14553 8619 14611 8625
rect 14553 8616 14565 8619
rect 14424 8588 14565 8616
rect 14424 8576 14430 8588
rect 14553 8585 14565 8588
rect 14599 8585 14611 8619
rect 14553 8579 14611 8585
rect 17770 8576 17776 8628
rect 17828 8576 17834 8628
rect 20070 8616 20076 8628
rect 18616 8588 20076 8616
rect 6181 8551 6239 8557
rect 6181 8548 6193 8551
rect 5920 8520 6193 8548
rect 6181 8517 6193 8520
rect 6227 8517 6239 8551
rect 6181 8511 6239 8517
rect 10870 8508 10876 8560
rect 10928 8508 10934 8560
rect 10962 8508 10968 8560
rect 11020 8548 11026 8560
rect 11885 8551 11943 8557
rect 11885 8548 11897 8551
rect 11020 8520 11897 8548
rect 11020 8508 11026 8520
rect 11885 8517 11897 8520
rect 11931 8517 11943 8551
rect 11885 8511 11943 8517
rect 13725 8551 13783 8557
rect 13725 8517 13737 8551
rect 13771 8548 13783 8551
rect 14642 8548 14648 8560
rect 13771 8520 14648 8548
rect 13771 8517 13783 8520
rect 13725 8511 13783 8517
rect 14642 8508 14648 8520
rect 14700 8508 14706 8560
rect 14921 8551 14979 8557
rect 14921 8517 14933 8551
rect 14967 8548 14979 8551
rect 15194 8548 15200 8560
rect 14967 8520 15200 8548
rect 14967 8517 14979 8520
rect 14921 8511 14979 8517
rect 15194 8508 15200 8520
rect 15252 8508 15258 8560
rect 6362 8440 6368 8492
rect 6420 8440 6426 8492
rect 9858 8480 9864 8492
rect 9048 8452 9864 8480
rect 6380 8412 6408 8440
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 6380 8384 6561 8412
rect 6549 8381 6561 8384
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 7926 8372 7932 8424
rect 7984 8372 7990 8424
rect 8110 8372 8116 8424
rect 8168 8372 8174 8424
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8478 8412 8484 8424
rect 8251 8384 8484 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 5074 8304 5080 8356
rect 5132 8344 5138 8356
rect 6365 8347 6423 8353
rect 6365 8344 6377 8347
rect 5132 8316 6377 8344
rect 5132 8304 5138 8316
rect 6365 8313 6377 8316
rect 6411 8313 6423 8347
rect 6365 8307 6423 8313
rect 7190 8304 7196 8356
rect 7248 8344 7254 8356
rect 8220 8344 8248 8375
rect 8478 8372 8484 8384
rect 8536 8372 8542 8424
rect 9048 8421 9076 8452
rect 9858 8440 9864 8452
rect 9916 8480 9922 8492
rect 10980 8480 11008 8508
rect 9916 8452 11008 8480
rect 9916 8440 9922 8452
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 14550 8480 14556 8492
rect 13044 8452 14556 8480
rect 13044 8440 13050 8452
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 10870 8372 10876 8424
rect 10928 8412 10934 8424
rect 11425 8415 11483 8421
rect 11425 8412 11437 8415
rect 10928 8384 11437 8412
rect 10928 8372 10934 8384
rect 11425 8381 11437 8384
rect 11471 8381 11483 8415
rect 11425 8375 11483 8381
rect 11514 8372 11520 8424
rect 11572 8412 11578 8424
rect 11609 8415 11667 8421
rect 11609 8412 11621 8415
rect 11572 8384 11621 8412
rect 11572 8372 11578 8384
rect 11609 8381 11621 8384
rect 11655 8412 11667 8415
rect 11790 8412 11796 8424
rect 11655 8384 11796 8412
rect 11655 8381 11667 8384
rect 11609 8375 11667 8381
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 13372 8421 13400 8452
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 16393 8483 16451 8489
rect 16393 8480 16405 8483
rect 16356 8452 16405 8480
rect 16356 8440 16362 8452
rect 16393 8449 16405 8452
rect 16439 8449 16451 8483
rect 16393 8443 16451 8449
rect 17402 8440 17408 8492
rect 17460 8480 17466 8492
rect 17460 8452 18092 8480
rect 17460 8440 17466 8452
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 11940 8384 12081 8412
rect 11940 8372 11946 8384
rect 12069 8381 12081 8384
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 13173 8415 13231 8421
rect 13173 8381 13185 8415
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8381 13415 8415
rect 13357 8375 13415 8381
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8412 14335 8415
rect 14323 8384 14780 8412
rect 14323 8381 14335 8384
rect 14277 8375 14335 8381
rect 7248 8316 8248 8344
rect 7248 8304 7254 8316
rect 8386 8304 8392 8356
rect 8444 8304 8450 8356
rect 8570 8304 8576 8356
rect 8628 8304 8634 8356
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 11146 8344 11152 8356
rect 10744 8316 11152 8344
rect 10744 8304 10750 8316
rect 11146 8304 11152 8316
rect 11204 8344 11210 8356
rect 11241 8347 11299 8353
rect 11241 8344 11253 8347
rect 11204 8316 11253 8344
rect 11204 8304 11210 8316
rect 11241 8313 11253 8316
rect 11287 8344 11299 8347
rect 12342 8344 12348 8356
rect 11287 8316 12348 8344
rect 11287 8313 11299 8316
rect 11241 8307 11299 8313
rect 12342 8304 12348 8316
rect 12400 8304 12406 8356
rect 13078 8304 13084 8356
rect 13136 8344 13142 8356
rect 13188 8344 13216 8375
rect 13722 8344 13728 8356
rect 13136 8316 13728 8344
rect 13136 8304 13142 8316
rect 13722 8304 13728 8316
rect 13780 8344 13786 8356
rect 14369 8347 14427 8353
rect 14369 8344 14381 8347
rect 13780 8316 14381 8344
rect 13780 8304 13786 8316
rect 14369 8313 14381 8316
rect 14415 8344 14427 8347
rect 14458 8344 14464 8356
rect 14415 8316 14464 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 14550 8304 14556 8356
rect 14608 8353 14614 8356
rect 14608 8347 14627 8353
rect 14615 8313 14627 8347
rect 14608 8307 14627 8313
rect 14608 8304 14614 8307
rect 14752 8288 14780 8384
rect 16482 8372 16488 8424
rect 16540 8412 16546 8424
rect 17420 8412 17448 8440
rect 16540 8384 17448 8412
rect 16540 8372 16546 8384
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 18064 8421 18092 8452
rect 17865 8415 17923 8421
rect 17865 8412 17877 8415
rect 17828 8384 17877 8412
rect 17828 8372 17834 8384
rect 17865 8381 17877 8384
rect 17911 8381 17923 8415
rect 17865 8375 17923 8381
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 18325 8415 18383 8421
rect 18325 8381 18337 8415
rect 18371 8412 18383 8415
rect 18616 8412 18644 8588
rect 20070 8576 20076 8588
rect 20128 8576 20134 8628
rect 20349 8619 20407 8625
rect 20349 8585 20361 8619
rect 20395 8616 20407 8619
rect 20898 8616 20904 8628
rect 20395 8588 20904 8616
rect 20395 8585 20407 8588
rect 20349 8579 20407 8585
rect 20364 8548 20392 8579
rect 20898 8576 20904 8588
rect 20956 8616 20962 8628
rect 21082 8616 21088 8628
rect 20956 8588 21088 8616
rect 20956 8576 20962 8588
rect 21082 8576 21088 8588
rect 21140 8616 21146 8628
rect 21361 8619 21419 8625
rect 21361 8616 21373 8619
rect 21140 8588 21373 8616
rect 21140 8576 21146 8588
rect 21361 8585 21373 8588
rect 21407 8585 21419 8619
rect 21361 8579 21419 8585
rect 22557 8619 22615 8625
rect 22557 8585 22569 8619
rect 22603 8585 22615 8619
rect 22557 8579 22615 8585
rect 20088 8520 20392 8548
rect 20717 8551 20775 8557
rect 18690 8440 18696 8492
rect 18748 8440 18754 8492
rect 18371 8384 18644 8412
rect 18371 8381 18383 8384
rect 18325 8375 18383 8381
rect 19242 8372 19248 8424
rect 19300 8412 19306 8424
rect 20088 8412 20116 8520
rect 20717 8517 20729 8551
rect 20763 8548 20775 8551
rect 22373 8551 22431 8557
rect 22373 8548 22385 8551
rect 20763 8520 22385 8548
rect 20763 8517 20775 8520
rect 20717 8511 20775 8517
rect 22373 8517 22385 8520
rect 22419 8517 22431 8551
rect 22373 8511 22431 8517
rect 20732 8412 20760 8511
rect 20806 8440 20812 8492
rect 20864 8480 20870 8492
rect 22572 8480 22600 8579
rect 20864 8452 22600 8480
rect 20864 8440 20870 8452
rect 19300 8384 20116 8412
rect 20180 8384 20760 8412
rect 20901 8415 20959 8421
rect 19300 8372 19306 8384
rect 15010 8304 15016 8356
rect 15068 8344 15074 8356
rect 16034 8347 16092 8353
rect 16034 8344 16046 8347
rect 15068 8316 16046 8344
rect 15068 8304 15074 8316
rect 16034 8313 16046 8316
rect 16080 8313 16092 8347
rect 16034 8307 16092 8313
rect 16660 8347 16718 8353
rect 16660 8313 16672 8347
rect 16706 8344 16718 8347
rect 16942 8344 16948 8356
rect 16706 8316 16948 8344
rect 16706 8313 16718 8316
rect 16660 8307 16718 8313
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 18509 8347 18567 8353
rect 18509 8313 18521 8347
rect 18555 8344 18567 8347
rect 18555 8316 18736 8344
rect 18555 8313 18567 8316
rect 18509 8307 18567 8313
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5905 8279 5963 8285
rect 5905 8276 5917 8279
rect 4948 8248 5917 8276
rect 4948 8236 4954 8248
rect 5905 8245 5917 8248
rect 5951 8276 5963 8279
rect 7558 8276 7564 8288
rect 5951 8248 7564 8276
rect 5951 8245 5963 8248
rect 5905 8239 5963 8245
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 7745 8279 7803 8285
rect 7745 8245 7757 8279
rect 7791 8276 7803 8279
rect 7834 8276 7840 8288
rect 7791 8248 7840 8276
rect 7791 8245 7803 8248
rect 7745 8239 7803 8245
rect 7834 8236 7840 8248
rect 7892 8236 7898 8288
rect 8757 8279 8815 8285
rect 8757 8245 8769 8279
rect 8803 8276 8815 8279
rect 8846 8276 8852 8288
rect 8803 8248 8852 8276
rect 8803 8245 8815 8248
rect 8757 8239 8815 8245
rect 8846 8236 8852 8248
rect 8904 8236 8910 8288
rect 8938 8236 8944 8288
rect 8996 8236 9002 8288
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 10594 8276 10600 8288
rect 9824 8248 10600 8276
rect 9824 8236 9830 8248
rect 10594 8236 10600 8248
rect 10652 8276 10658 8288
rect 11054 8285 11060 8288
rect 11031 8279 11060 8285
rect 11031 8276 11043 8279
rect 10652 8248 11043 8276
rect 10652 8236 10658 8248
rect 11031 8245 11043 8248
rect 11112 8276 11118 8288
rect 11606 8276 11612 8288
rect 11112 8248 11612 8276
rect 11031 8239 11060 8245
rect 11054 8236 11060 8239
rect 11112 8236 11118 8248
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 11790 8236 11796 8288
rect 11848 8236 11854 8288
rect 13170 8236 13176 8288
rect 13228 8236 13234 8288
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 13909 8279 13967 8285
rect 13909 8276 13921 8279
rect 13504 8248 13921 8276
rect 13504 8236 13510 8248
rect 13909 8245 13921 8248
rect 13955 8276 13967 8279
rect 14274 8276 14280 8288
rect 13955 8248 14280 8276
rect 13955 8245 13967 8248
rect 13909 8239 13967 8245
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 14734 8236 14740 8288
rect 14792 8236 14798 8288
rect 17954 8236 17960 8288
rect 18012 8236 18018 8288
rect 18138 8236 18144 8288
rect 18196 8236 18202 8288
rect 18708 8276 18736 8316
rect 18782 8304 18788 8356
rect 18840 8344 18846 8356
rect 18938 8347 18996 8353
rect 18938 8344 18950 8347
rect 18840 8316 18950 8344
rect 18840 8304 18846 8316
rect 18938 8313 18950 8316
rect 18984 8313 18996 8347
rect 19426 8344 19432 8356
rect 18938 8307 18996 8313
rect 19076 8316 19432 8344
rect 19076 8276 19104 8316
rect 19426 8304 19432 8316
rect 19484 8344 19490 8356
rect 20180 8344 20208 8384
rect 20901 8381 20913 8415
rect 20947 8412 20959 8415
rect 20990 8412 20996 8424
rect 20947 8384 20996 8412
rect 20947 8381 20959 8384
rect 20901 8375 20959 8381
rect 20990 8372 20996 8384
rect 21048 8372 21054 8424
rect 21085 8415 21143 8421
rect 21085 8381 21097 8415
rect 21131 8412 21143 8415
rect 21634 8412 21640 8424
rect 21131 8384 21640 8412
rect 21131 8381 21143 8384
rect 21085 8375 21143 8381
rect 21634 8372 21640 8384
rect 21692 8412 21698 8424
rect 22020 8421 22048 8452
rect 21729 8415 21787 8421
rect 21729 8412 21741 8415
rect 21692 8384 21741 8412
rect 21692 8372 21698 8384
rect 21729 8381 21741 8384
rect 21775 8381 21787 8415
rect 21729 8375 21787 8381
rect 22005 8415 22063 8421
rect 22005 8381 22017 8415
rect 22051 8381 22063 8415
rect 22005 8375 22063 8381
rect 22281 8415 22339 8421
rect 22281 8381 22293 8415
rect 22327 8381 22339 8415
rect 22281 8375 22339 8381
rect 19484 8316 20208 8344
rect 20349 8347 20407 8353
rect 19484 8304 19490 8316
rect 20349 8313 20361 8347
rect 20395 8344 20407 8347
rect 21821 8347 21879 8353
rect 21821 8344 21833 8347
rect 20395 8316 21833 8344
rect 20395 8313 20407 8316
rect 20349 8307 20407 8313
rect 21821 8313 21833 8316
rect 21867 8313 21879 8347
rect 21821 8307 21879 8313
rect 21910 8304 21916 8356
rect 21968 8344 21974 8356
rect 22189 8347 22247 8353
rect 22189 8344 22201 8347
rect 21968 8316 22201 8344
rect 21968 8304 21974 8316
rect 22189 8313 22201 8316
rect 22235 8313 22247 8347
rect 22189 8307 22247 8313
rect 18708 8248 19104 8276
rect 20162 8236 20168 8288
rect 20220 8236 20226 8288
rect 20993 8279 21051 8285
rect 20993 8245 21005 8279
rect 21039 8276 21051 8279
rect 21082 8276 21088 8288
rect 21039 8248 21088 8276
rect 21039 8245 21051 8248
rect 20993 8239 21051 8245
rect 21082 8236 21088 8248
rect 21140 8236 21146 8288
rect 21174 8236 21180 8288
rect 21232 8236 21238 8288
rect 21266 8236 21272 8288
rect 21324 8276 21330 8288
rect 21361 8279 21419 8285
rect 21361 8276 21373 8279
rect 21324 8248 21373 8276
rect 21324 8236 21330 8248
rect 21361 8245 21373 8248
rect 21407 8245 21419 8279
rect 21361 8239 21419 8245
rect 21634 8236 21640 8288
rect 21692 8276 21698 8288
rect 22296 8276 22324 8375
rect 22646 8304 22652 8356
rect 22704 8344 22710 8356
rect 22741 8347 22799 8353
rect 22741 8344 22753 8347
rect 22704 8316 22753 8344
rect 22704 8304 22710 8316
rect 22741 8313 22753 8316
rect 22787 8313 22799 8347
rect 22741 8307 22799 8313
rect 22541 8279 22599 8285
rect 22541 8276 22553 8279
rect 21692 8248 22553 8276
rect 21692 8236 21698 8248
rect 22541 8245 22553 8248
rect 22587 8245 22599 8279
rect 22541 8239 22599 8245
rect 552 8186 23368 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 23368 8186
rect 552 8112 23368 8134
rect 7190 8072 7196 8084
rect 7248 8081 7254 8084
rect 7248 8075 7272 8081
rect 6748 8044 7196 8072
rect 4246 7964 4252 8016
rect 4304 7964 4310 8016
rect 4709 8007 4767 8013
rect 4709 7973 4721 8007
rect 4755 7973 4767 8007
rect 4709 7967 4767 7973
rect 4925 8007 4983 8013
rect 4925 7973 4937 8007
rect 4971 8004 4983 8007
rect 5626 8004 5632 8016
rect 4971 7976 5632 8004
rect 4971 7973 4983 7976
rect 4925 7967 4983 7973
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 4724 7936 4752 7967
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 3568 7908 4752 7936
rect 3568 7896 3574 7908
rect 5718 7896 5724 7948
rect 5776 7936 5782 7948
rect 6748 7945 6776 8044
rect 7190 8032 7196 8044
rect 7260 8041 7272 8075
rect 7248 8035 7272 8041
rect 7377 8075 7435 8081
rect 7377 8041 7389 8075
rect 7423 8072 7435 8075
rect 8386 8072 8392 8084
rect 7423 8044 8392 8072
rect 7423 8041 7435 8044
rect 7377 8035 7435 8041
rect 7248 8032 7254 8035
rect 7009 8007 7067 8013
rect 7009 7973 7021 8007
rect 7055 7973 7067 8007
rect 7009 7967 7067 7973
rect 6733 7939 6791 7945
rect 6733 7936 6745 7939
rect 5776 7908 6745 7936
rect 5776 7896 5782 7908
rect 6733 7905 6745 7908
rect 6779 7905 6791 7939
rect 6733 7899 6791 7905
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7936 6975 7939
rect 7024 7936 7052 7967
rect 7484 7945 7512 8044
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8478 8032 8484 8084
rect 8536 8032 8542 8084
rect 10686 8032 10692 8084
rect 10744 8032 10750 8084
rect 11330 8032 11336 8084
rect 11388 8072 11394 8084
rect 11425 8075 11483 8081
rect 11425 8072 11437 8075
rect 11388 8044 11437 8072
rect 11388 8032 11394 8044
rect 11425 8041 11437 8044
rect 11471 8041 11483 8075
rect 11425 8035 11483 8041
rect 11514 8032 11520 8084
rect 11572 8032 11578 8084
rect 13078 8032 13084 8084
rect 13136 8032 13142 8084
rect 13449 8075 13507 8081
rect 13449 8041 13461 8075
rect 13495 8072 13507 8075
rect 13906 8072 13912 8084
rect 13495 8044 13912 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14332 8044 14964 8072
rect 14332 8032 14338 8044
rect 7558 7964 7564 8016
rect 7616 8004 7622 8016
rect 7837 8007 7895 8013
rect 7837 8004 7849 8007
rect 7616 7976 7849 8004
rect 7616 7964 7622 7976
rect 7837 7973 7849 7976
rect 7883 7973 7895 8007
rect 7837 7967 7895 7973
rect 6963 7908 7052 7936
rect 6963 7905 6975 7908
rect 6917 7899 6975 7905
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 5442 7868 5448 7880
rect 4663 7840 5448 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 7024 7868 7052 7908
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7905 7527 7939
rect 7852 7936 7880 7967
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 8297 8007 8355 8013
rect 8297 8004 8309 8007
rect 7984 7976 8309 8004
rect 7984 7964 7990 7976
rect 8297 7973 8309 7976
rect 8343 7973 8355 8007
rect 8297 7967 8355 7973
rect 8941 8007 8999 8013
rect 8941 7973 8953 8007
rect 8987 8004 8999 8007
rect 9861 8007 9919 8013
rect 9861 8004 9873 8007
rect 8987 7976 9873 8004
rect 8987 7973 8999 7976
rect 8941 7967 8999 7973
rect 9861 7973 9873 7976
rect 9907 8004 9919 8007
rect 9950 8004 9956 8016
rect 9907 7976 9956 8004
rect 9907 7973 9919 7976
rect 9861 7967 9919 7973
rect 9950 7964 9956 7976
rect 10008 7964 10014 8016
rect 10077 8007 10135 8013
rect 10077 7973 10089 8007
rect 10123 8004 10135 8007
rect 10318 8004 10324 8016
rect 10123 7976 10324 8004
rect 10123 7973 10135 7976
rect 10077 7967 10135 7973
rect 10318 7964 10324 7976
rect 10376 7964 10382 8016
rect 10765 7961 10823 7967
rect 11698 7964 11704 8016
rect 11756 8004 11762 8016
rect 12253 8007 12311 8013
rect 12253 8004 12265 8007
rect 11756 7976 12265 8004
rect 11756 7964 11762 7976
rect 12253 7973 12265 7976
rect 12299 8004 12311 8007
rect 12529 8007 12587 8013
rect 12529 8004 12541 8007
rect 12299 7976 12541 8004
rect 12299 7973 12311 7976
rect 12253 7967 12311 7973
rect 12529 7973 12541 7976
rect 12575 7973 12587 8007
rect 12529 7967 12587 7973
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 12768 7976 14504 8004
rect 12768 7964 12774 7976
rect 10765 7958 10777 7961
rect 10612 7948 10777 7958
rect 8018 7936 8024 7948
rect 7852 7908 8024 7936
rect 7469 7899 7527 7905
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 8110 7896 8116 7948
rect 8168 7896 8174 7948
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 7190 7868 7196 7880
rect 7024 7840 7196 7868
rect 7190 7828 7196 7840
rect 7248 7868 7254 7880
rect 8128 7868 8156 7896
rect 7248 7840 8156 7868
rect 8404 7868 8432 7899
rect 10502 7896 10508 7948
rect 10560 7896 10566 7948
rect 10594 7896 10600 7948
rect 10652 7930 10777 7948
rect 10652 7896 10658 7930
rect 10765 7927 10777 7930
rect 10811 7927 10823 7961
rect 10765 7921 10823 7927
rect 10965 7937 11023 7943
rect 10965 7903 10977 7937
rect 11011 7903 11023 7937
rect 10965 7897 11023 7903
rect 8570 7868 8576 7880
rect 8404 7840 8576 7868
rect 7248 7828 7254 7840
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 10980 7868 11008 7897
rect 11054 7896 11060 7948
rect 11112 7936 11118 7948
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 11112 7908 11161 7936
rect 11112 7896 11118 7908
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 11149 7899 11207 7905
rect 11238 7896 11244 7948
rect 11296 7896 11302 7948
rect 11606 7896 11612 7948
rect 11664 7896 11670 7948
rect 12986 7896 12992 7948
rect 13044 7896 13050 7948
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7936 13323 7939
rect 14366 7936 14372 7948
rect 13311 7908 14372 7936
rect 13311 7905 13323 7908
rect 13265 7899 13323 7905
rect 11793 7871 11851 7877
rect 10980 7840 11100 7868
rect 7558 7800 7564 7812
rect 7208 7772 7564 7800
rect 4062 7692 4068 7744
rect 4120 7692 4126 7744
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 4212 7704 4261 7732
rect 4212 7692 4218 7704
rect 4249 7701 4261 7704
rect 4295 7732 4307 7735
rect 4890 7732 4896 7744
rect 4295 7704 4896 7732
rect 4295 7701 4307 7704
rect 4249 7695 4307 7701
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5074 7692 5080 7744
rect 5132 7692 5138 7744
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 7208 7741 7236 7772
rect 7558 7760 7564 7772
rect 7616 7800 7622 7812
rect 7926 7800 7932 7812
rect 7616 7772 7932 7800
rect 7616 7760 7622 7772
rect 7926 7760 7932 7772
rect 7984 7760 7990 7812
rect 8665 7803 8723 7809
rect 8665 7769 8677 7803
rect 8711 7800 8723 7803
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 8711 7772 9321 7800
rect 8711 7769 8723 7772
rect 8665 7763 8723 7769
rect 9309 7769 9321 7772
rect 9355 7800 9367 7803
rect 9766 7800 9772 7812
rect 9355 7772 9772 7800
rect 9355 7769 9367 7772
rect 9309 7763 9367 7769
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 11072 7800 11100 7840
rect 11793 7837 11805 7871
rect 11839 7868 11851 7871
rect 11885 7871 11943 7877
rect 11885 7868 11897 7871
rect 11839 7840 11897 7868
rect 11839 7837 11851 7840
rect 11793 7831 11851 7837
rect 11885 7837 11897 7840
rect 11931 7868 11943 7871
rect 13004 7868 13032 7896
rect 11931 7840 13032 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 11146 7800 11152 7812
rect 10060 7772 10548 7800
rect 11072 7772 11152 7800
rect 6825 7735 6883 7741
rect 6825 7732 6837 7735
rect 6604 7704 6837 7732
rect 6604 7692 6610 7704
rect 6825 7701 6837 7704
rect 6871 7701 6883 7735
rect 6825 7695 6883 7701
rect 7193 7735 7251 7741
rect 7193 7701 7205 7735
rect 7239 7701 7251 7735
rect 7193 7695 7251 7701
rect 7834 7692 7840 7744
rect 7892 7692 7898 7744
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 8386 7732 8392 7744
rect 8067 7704 8392 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 8754 7692 8760 7744
rect 8812 7692 8818 7744
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 10060 7741 10088 7772
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8904 7704 8953 7732
rect 8904 7692 8910 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 8941 7695 8999 7701
rect 10045 7735 10103 7741
rect 10045 7701 10057 7735
rect 10091 7701 10103 7735
rect 10045 7695 10103 7701
rect 10226 7692 10232 7744
rect 10284 7692 10290 7744
rect 10321 7735 10379 7741
rect 10321 7701 10333 7735
rect 10367 7732 10379 7735
rect 10410 7732 10416 7744
rect 10367 7704 10416 7732
rect 10367 7701 10379 7704
rect 10321 7695 10379 7701
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 10520 7732 10548 7772
rect 11146 7760 11152 7772
rect 11204 7760 11210 7812
rect 13280 7800 13308 7899
rect 14366 7896 14372 7908
rect 14424 7896 14430 7948
rect 14476 7936 14504 7976
rect 14642 7964 14648 8016
rect 14700 8013 14706 8016
rect 14700 8004 14712 8013
rect 14936 8004 14964 8044
rect 15010 8032 15016 8084
rect 15068 8032 15074 8084
rect 16666 8072 16672 8084
rect 15212 8044 16672 8072
rect 15212 8013 15240 8044
rect 16666 8032 16672 8044
rect 16724 8072 16730 8084
rect 16724 8044 17356 8072
rect 16724 8032 16730 8044
rect 15197 8007 15255 8013
rect 15197 8004 15209 8007
rect 14700 7976 14745 8004
rect 14936 7976 15209 8004
rect 14700 7967 14712 7976
rect 15197 7973 15209 7976
rect 15243 7973 15255 8007
rect 15197 7967 15255 7973
rect 14700 7964 14706 7967
rect 16482 7964 16488 8016
rect 16540 7964 16546 8016
rect 17328 8013 17356 8044
rect 18782 8032 18788 8084
rect 18840 8032 18846 8084
rect 19518 8032 19524 8084
rect 19576 8032 19582 8084
rect 19886 8032 19892 8084
rect 19944 8032 19950 8084
rect 20806 8032 20812 8084
rect 20864 8072 20870 8084
rect 21085 8075 21143 8081
rect 21085 8072 21097 8075
rect 20864 8044 21097 8072
rect 20864 8032 20870 8044
rect 21085 8041 21097 8044
rect 21131 8041 21143 8075
rect 21085 8035 21143 8041
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 22646 8072 22652 8084
rect 21968 8044 22652 8072
rect 21968 8032 21974 8044
rect 22646 8032 22652 8044
rect 22704 8032 22710 8084
rect 16853 8007 16911 8013
rect 16853 7973 16865 8007
rect 16899 8004 16911 8007
rect 17097 8007 17155 8013
rect 17097 8004 17109 8007
rect 16899 7976 17109 8004
rect 16899 7973 16911 7976
rect 16853 7967 16911 7973
rect 17097 7973 17109 7976
rect 17143 7973 17155 8007
rect 17097 7967 17155 7973
rect 17313 8007 17371 8013
rect 17313 7973 17325 8007
rect 17359 7973 17371 8007
rect 17313 7967 17371 7973
rect 18138 7964 18144 8016
rect 18196 8004 18202 8016
rect 18969 8007 19027 8013
rect 18969 8004 18981 8007
rect 18196 7976 18981 8004
rect 18196 7964 18202 7976
rect 18969 7973 18981 7976
rect 19015 7973 19027 8007
rect 18969 7967 19027 7973
rect 14476 7908 14872 7936
rect 14844 7868 14872 7908
rect 14918 7896 14924 7948
rect 14976 7896 14982 7948
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7936 16727 7939
rect 17770 7936 17776 7948
rect 16715 7908 17776 7936
rect 16715 7905 16727 7908
rect 16669 7899 16727 7905
rect 17770 7896 17776 7908
rect 17828 7896 17834 7948
rect 19337 7939 19395 7945
rect 19337 7905 19349 7939
rect 19383 7936 19395 7939
rect 19429 7939 19487 7945
rect 19429 7936 19441 7939
rect 19383 7908 19441 7936
rect 19383 7905 19395 7908
rect 19337 7899 19395 7905
rect 19429 7905 19441 7908
rect 19475 7936 19487 7939
rect 19518 7936 19524 7948
rect 19475 7908 19524 7936
rect 19475 7905 19487 7908
rect 19429 7899 19487 7905
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 19613 7939 19671 7945
rect 19613 7905 19625 7939
rect 19659 7936 19671 7939
rect 19904 7936 19932 8032
rect 19972 8007 20030 8013
rect 19972 7973 19984 8007
rect 20018 8004 20030 8007
rect 20162 8004 20168 8016
rect 20018 7976 20168 8004
rect 20018 7973 20030 7976
rect 19972 7967 20030 7973
rect 20162 7964 20168 7976
rect 20220 7964 20226 8016
rect 20990 7964 20996 8016
rect 21048 8004 21054 8016
rect 21358 8004 21364 8016
rect 21048 7976 21364 8004
rect 21048 7964 21054 7976
rect 21358 7964 21364 7976
rect 21416 8004 21422 8016
rect 21928 8004 21956 8032
rect 21416 7976 21956 8004
rect 21416 7964 21422 7976
rect 22002 7964 22008 8016
rect 22060 8004 22066 8016
rect 22741 8007 22799 8013
rect 22741 8004 22753 8007
rect 22060 7976 22753 8004
rect 22060 7964 22066 7976
rect 22741 7973 22753 7976
rect 22787 7973 22799 8007
rect 22741 7967 22799 7973
rect 21542 7945 21548 7948
rect 19659 7908 19932 7936
rect 19659 7905 19671 7908
rect 19613 7899 19671 7905
rect 21536 7899 21548 7945
rect 21542 7896 21548 7899
rect 21600 7896 21606 7948
rect 21818 7896 21824 7948
rect 21876 7936 21882 7948
rect 22925 7939 22983 7945
rect 22925 7936 22937 7939
rect 21876 7908 22937 7936
rect 21876 7896 21882 7908
rect 22925 7905 22937 7908
rect 22971 7905 22983 7939
rect 22925 7899 22983 7905
rect 14844 7840 19334 7868
rect 13541 7803 13599 7809
rect 13541 7800 13553 7803
rect 13280 7772 13553 7800
rect 13541 7769 13553 7772
rect 13587 7769 13599 7803
rect 13541 7763 13599 7769
rect 15565 7803 15623 7809
rect 15565 7769 15577 7803
rect 15611 7800 15623 7803
rect 16482 7800 16488 7812
rect 15611 7772 16488 7800
rect 15611 7769 15623 7772
rect 15565 7763 15623 7769
rect 16482 7760 16488 7772
rect 16540 7760 16546 7812
rect 16942 7760 16948 7812
rect 17000 7760 17006 7812
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10520 7704 11069 7732
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 11790 7692 11796 7744
rect 11848 7732 11854 7744
rect 12253 7735 12311 7741
rect 12253 7732 12265 7735
rect 11848 7704 12265 7732
rect 11848 7692 11854 7704
rect 12253 7701 12265 7704
rect 12299 7701 12311 7735
rect 12253 7695 12311 7701
rect 12434 7692 12440 7744
rect 12492 7692 12498 7744
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 14918 7732 14924 7744
rect 13412 7704 14924 7732
rect 13412 7692 13418 7704
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 15197 7735 15255 7741
rect 15197 7701 15209 7735
rect 15243 7732 15255 7735
rect 15378 7732 15384 7744
rect 15243 7704 15384 7732
rect 15243 7701 15255 7704
rect 15197 7695 15255 7701
rect 15378 7692 15384 7704
rect 15436 7692 15442 7744
rect 17129 7735 17187 7741
rect 17129 7701 17141 7735
rect 17175 7732 17187 7735
rect 17954 7732 17960 7744
rect 17175 7704 17960 7732
rect 17175 7701 17187 7704
rect 17129 7695 17187 7701
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18969 7735 19027 7741
rect 18969 7701 18981 7735
rect 19015 7732 19027 7735
rect 19150 7732 19156 7744
rect 19015 7704 19156 7732
rect 19015 7701 19027 7704
rect 18969 7695 19027 7701
rect 19150 7692 19156 7704
rect 19208 7692 19214 7744
rect 19306 7732 19334 7840
rect 19702 7828 19708 7880
rect 19760 7828 19766 7880
rect 21269 7871 21327 7877
rect 21269 7837 21281 7871
rect 21315 7837 21327 7871
rect 21269 7831 21327 7837
rect 20714 7732 20720 7744
rect 19306 7704 20720 7732
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 21284 7732 21312 7831
rect 22002 7732 22008 7744
rect 21284 7704 22008 7732
rect 22002 7692 22008 7704
rect 22060 7692 22066 7744
rect 552 7642 23368 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 23368 7642
rect 552 7568 23368 7590
rect 3510 7488 3516 7540
rect 3568 7488 3574 7540
rect 3602 7488 3608 7540
rect 3660 7528 3666 7540
rect 3881 7531 3939 7537
rect 3881 7528 3893 7531
rect 3660 7500 3893 7528
rect 3660 7488 3666 7500
rect 3881 7497 3893 7500
rect 3927 7528 3939 7531
rect 4154 7528 4160 7540
rect 3927 7500 4160 7528
rect 3927 7497 3939 7500
rect 3881 7491 3939 7497
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 5626 7488 5632 7540
rect 5684 7488 5690 7540
rect 6546 7488 6552 7540
rect 6604 7488 6610 7540
rect 8110 7488 8116 7540
rect 8168 7528 8174 7540
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 8168 7500 8217 7528
rect 8168 7488 8174 7500
rect 8205 7497 8217 7500
rect 8251 7497 8263 7531
rect 8205 7491 8263 7497
rect 8570 7488 8576 7540
rect 8628 7528 8634 7540
rect 9769 7531 9827 7537
rect 9769 7528 9781 7531
rect 8628 7500 9781 7528
rect 8628 7488 8634 7500
rect 9769 7497 9781 7500
rect 9815 7497 9827 7531
rect 9769 7491 9827 7497
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 11054 7528 11060 7540
rect 10284 7500 11060 7528
rect 10284 7488 10290 7500
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 11238 7488 11244 7540
rect 11296 7488 11302 7540
rect 11333 7531 11391 7537
rect 11333 7497 11345 7531
rect 11379 7528 11391 7531
rect 11514 7528 11520 7540
rect 11379 7500 11520 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 13170 7488 13176 7540
rect 13228 7488 13234 7540
rect 13538 7488 13544 7540
rect 13596 7528 13602 7540
rect 14458 7528 14464 7540
rect 13596 7500 14464 7528
rect 13596 7488 13602 7500
rect 14458 7488 14464 7500
rect 14516 7528 14522 7540
rect 14921 7531 14979 7537
rect 14921 7528 14933 7531
rect 14516 7500 14933 7528
rect 14516 7488 14522 7500
rect 14921 7497 14933 7500
rect 14967 7497 14979 7531
rect 14921 7491 14979 7497
rect 15378 7488 15384 7540
rect 15436 7488 15442 7540
rect 19245 7531 19303 7537
rect 19245 7497 19257 7531
rect 19291 7528 19303 7531
rect 19518 7528 19524 7540
rect 19291 7500 19524 7528
rect 19291 7497 19303 7500
rect 19245 7491 19303 7497
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 21542 7488 21548 7540
rect 21600 7528 21606 7540
rect 21637 7531 21695 7537
rect 21637 7528 21649 7531
rect 21600 7500 21649 7528
rect 21600 7488 21606 7500
rect 21637 7497 21649 7500
rect 21683 7497 21695 7531
rect 21637 7491 21695 7497
rect 21818 7488 21824 7540
rect 21876 7488 21882 7540
rect 4062 7420 4068 7472
rect 4120 7420 4126 7472
rect 6733 7463 6791 7469
rect 6733 7429 6745 7463
rect 6779 7429 6791 7463
rect 13446 7460 13452 7472
rect 6733 7423 6791 7429
rect 13004 7432 13452 7460
rect 3326 7352 3332 7404
rect 3384 7392 3390 7404
rect 4080 7392 4108 7420
rect 3384 7364 3648 7392
rect 4080 7364 4292 7392
rect 3384 7352 3390 7364
rect 3234 7284 3240 7336
rect 3292 7324 3298 7336
rect 3620 7333 3648 7364
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3292 7296 3433 7324
rect 3292 7284 3298 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7293 3663 7327
rect 3605 7287 3663 7293
rect 4062 7284 4068 7336
rect 4120 7284 4126 7336
rect 4157 7327 4215 7333
rect 4157 7293 4169 7327
rect 4203 7293 4215 7327
rect 4264 7324 4292 7364
rect 4413 7327 4471 7333
rect 4413 7324 4425 7327
rect 4264 7296 4425 7324
rect 4157 7287 4215 7293
rect 4413 7293 4425 7296
rect 4459 7293 4471 7327
rect 4413 7287 4471 7293
rect 3697 7259 3755 7265
rect 3697 7256 3709 7259
rect 3436 7228 3709 7256
rect 3436 7200 3464 7228
rect 3697 7225 3709 7228
rect 3743 7225 3755 7259
rect 3697 7219 3755 7225
rect 3913 7259 3971 7265
rect 3913 7225 3925 7259
rect 3959 7256 3971 7259
rect 4080 7256 4108 7284
rect 3959 7228 4108 7256
rect 4172 7256 4200 7287
rect 4706 7256 4712 7268
rect 4172 7228 4712 7256
rect 3959 7225 3971 7228
rect 3913 7219 3971 7225
rect 4706 7216 4712 7228
rect 4764 7256 4770 7268
rect 5718 7256 5724 7268
rect 4764 7228 5724 7256
rect 4764 7216 4770 7228
rect 5718 7216 5724 7228
rect 5776 7216 5782 7268
rect 5810 7216 5816 7268
rect 5868 7216 5874 7268
rect 5994 7216 6000 7268
rect 6052 7216 6058 7268
rect 6365 7259 6423 7265
rect 6365 7225 6377 7259
rect 6411 7256 6423 7259
rect 6748 7256 6776 7423
rect 9858 7352 9864 7404
rect 9916 7352 9922 7404
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 6880 7296 8401 7324
rect 6880 7284 6886 7296
rect 8389 7293 8401 7296
rect 8435 7324 8447 7327
rect 8938 7324 8944 7336
rect 8435 7296 8944 7324
rect 8435 7293 8447 7296
rect 8389 7287 8447 7293
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 12434 7284 12440 7336
rect 12492 7333 12498 7336
rect 12492 7324 12504 7333
rect 12713 7327 12771 7333
rect 12492 7296 12537 7324
rect 12492 7287 12504 7296
rect 12713 7293 12725 7327
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12492 7284 12498 7287
rect 7070 7259 7128 7265
rect 7070 7256 7082 7259
rect 6411 7228 6684 7256
rect 6748 7228 7082 7256
rect 6411 7225 6423 7228
rect 6365 7219 6423 7225
rect 3418 7148 3424 7200
rect 3476 7148 3482 7200
rect 4065 7191 4123 7197
rect 4065 7157 4077 7191
rect 4111 7188 4123 7191
rect 4154 7188 4160 7200
rect 4111 7160 4160 7188
rect 4111 7157 4123 7160
rect 4065 7151 4123 7157
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 5534 7148 5540 7200
rect 5592 7148 5598 7200
rect 6546 7148 6552 7200
rect 6604 7197 6610 7200
rect 6604 7191 6623 7197
rect 6611 7157 6623 7191
rect 6656 7188 6684 7228
rect 7070 7225 7082 7228
rect 7116 7225 7128 7259
rect 7070 7219 7128 7225
rect 8656 7259 8714 7265
rect 8656 7225 8668 7259
rect 8702 7256 8714 7259
rect 8754 7256 8760 7268
rect 8702 7228 8760 7256
rect 8702 7225 8714 7228
rect 8656 7219 8714 7225
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 10128 7259 10186 7265
rect 10128 7225 10140 7259
rect 10174 7256 10186 7259
rect 10226 7256 10232 7268
rect 10174 7228 10232 7256
rect 10174 7225 10186 7228
rect 10128 7219 10186 7225
rect 10226 7216 10232 7228
rect 10284 7216 10290 7268
rect 10962 7216 10968 7268
rect 11020 7256 11026 7268
rect 12728 7256 12756 7287
rect 13004 7265 13032 7432
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 19613 7395 19671 7401
rect 13096 7364 13676 7392
rect 11020 7228 12756 7256
rect 12989 7259 13047 7265
rect 11020 7216 11026 7228
rect 12989 7225 13001 7259
rect 13035 7225 13047 7259
rect 12989 7219 13047 7225
rect 8018 7188 8024 7200
rect 6656 7160 8024 7188
rect 6604 7151 6623 7157
rect 6604 7148 6610 7151
rect 8018 7148 8024 7160
rect 8076 7188 8082 7200
rect 11698 7188 11704 7200
rect 8076 7160 11704 7188
rect 8076 7148 8082 7160
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 11882 7148 11888 7200
rect 11940 7188 11946 7200
rect 13096 7188 13124 7364
rect 13354 7284 13360 7336
rect 13412 7324 13418 7336
rect 13541 7327 13599 7333
rect 13541 7324 13553 7327
rect 13412 7296 13553 7324
rect 13412 7284 13418 7296
rect 13541 7293 13553 7296
rect 13587 7293 13599 7327
rect 13648 7324 13676 7364
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 20070 7392 20076 7404
rect 19659 7364 20076 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 21634 7392 21640 7404
rect 21284 7364 21640 7392
rect 13648 7296 14688 7324
rect 13541 7287 13599 7293
rect 13786 7259 13844 7265
rect 13786 7256 13798 7259
rect 13648 7228 13798 7256
rect 11940 7160 13124 7188
rect 11940 7148 11946 7160
rect 13170 7148 13176 7200
rect 13228 7197 13234 7200
rect 13228 7191 13247 7197
rect 13235 7157 13247 7191
rect 13228 7151 13247 7157
rect 13357 7191 13415 7197
rect 13357 7157 13369 7191
rect 13403 7188 13415 7191
rect 13648 7188 13676 7228
rect 13786 7225 13798 7228
rect 13832 7225 13844 7259
rect 14660 7256 14688 7296
rect 14734 7284 14740 7336
rect 14792 7324 14798 7336
rect 15013 7327 15071 7333
rect 15013 7324 15025 7327
rect 14792 7296 15025 7324
rect 14792 7284 14798 7296
rect 15013 7293 15025 7296
rect 15059 7293 15071 7327
rect 15013 7287 15071 7293
rect 15194 7284 15200 7336
rect 15252 7284 15258 7336
rect 19426 7284 19432 7336
rect 19484 7284 19490 7336
rect 20898 7284 20904 7336
rect 20956 7324 20962 7336
rect 20993 7327 21051 7333
rect 20993 7324 21005 7327
rect 20956 7296 21005 7324
rect 20956 7284 20962 7296
rect 20993 7293 21005 7296
rect 21039 7293 21051 7327
rect 20993 7287 21051 7293
rect 21082 7284 21088 7336
rect 21140 7324 21146 7336
rect 21284 7333 21312 7364
rect 21634 7352 21640 7364
rect 21692 7352 21698 7404
rect 21177 7327 21235 7333
rect 21177 7324 21189 7327
rect 21140 7296 21189 7324
rect 21140 7284 21146 7296
rect 21177 7293 21189 7296
rect 21223 7293 21235 7327
rect 21177 7287 21235 7293
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7293 21327 7327
rect 21269 7287 21327 7293
rect 21358 7284 21364 7336
rect 21416 7284 21422 7336
rect 22738 7324 22744 7336
rect 22066 7296 22744 7324
rect 21913 7259 21971 7265
rect 21913 7256 21925 7259
rect 14660 7228 21925 7256
rect 13786 7219 13844 7225
rect 21913 7225 21925 7228
rect 21959 7256 21971 7259
rect 22066 7256 22094 7296
rect 22738 7284 22744 7296
rect 22796 7284 22802 7336
rect 21959 7228 22094 7256
rect 21959 7225 21971 7228
rect 21913 7219 21971 7225
rect 13403 7160 13676 7188
rect 13403 7157 13415 7160
rect 13357 7151 13415 7157
rect 13228 7148 13234 7151
rect 552 7098 23368 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 23368 7098
rect 552 7024 23368 7046
rect 4157 6987 4215 6993
rect 4157 6953 4169 6987
rect 4203 6984 4215 6987
rect 4246 6984 4252 6996
rect 4203 6956 4252 6984
rect 4203 6953 4215 6956
rect 4157 6947 4215 6953
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 5629 6987 5687 6993
rect 5629 6984 5641 6987
rect 5460 6956 5641 6984
rect 3234 6876 3240 6928
rect 3292 6916 3298 6928
rect 3786 6916 3792 6928
rect 3292 6888 3792 6916
rect 3292 6876 3298 6888
rect 3786 6876 3792 6888
rect 3844 6876 3850 6928
rect 4080 6888 4660 6916
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 3881 6851 3939 6857
rect 3881 6848 3893 6851
rect 3384 6820 3893 6848
rect 3384 6808 3390 6820
rect 3881 6817 3893 6820
rect 3927 6817 3939 6851
rect 3881 6811 3939 6817
rect 3973 6851 4031 6857
rect 3973 6817 3985 6851
rect 4019 6848 4031 6851
rect 4080 6848 4108 6888
rect 4019 6820 4108 6848
rect 4019 6817 4031 6820
rect 3973 6811 4031 6817
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6780 3111 6783
rect 3234 6780 3240 6792
rect 3099 6752 3240 6780
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3697 6783 3755 6789
rect 3697 6749 3709 6783
rect 3743 6749 3755 6783
rect 3697 6743 3755 6749
rect 3421 6715 3479 6721
rect 3421 6681 3433 6715
rect 3467 6712 3479 6715
rect 3602 6712 3608 6724
rect 3467 6684 3608 6712
rect 3467 6681 3479 6684
rect 3421 6675 3479 6681
rect 3602 6672 3608 6684
rect 3660 6672 3666 6724
rect 3510 6604 3516 6656
rect 3568 6604 3574 6656
rect 3712 6644 3740 6743
rect 3786 6740 3792 6792
rect 3844 6740 3850 6792
rect 4080 6712 4108 6820
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 4505 6851 4563 6857
rect 4505 6848 4517 6851
rect 4212 6820 4517 6848
rect 4212 6808 4218 6820
rect 4505 6817 4517 6820
rect 4551 6817 4563 6851
rect 4632 6848 4660 6888
rect 5460 6848 5488 6956
rect 5629 6953 5641 6956
rect 5675 6984 5687 6987
rect 6181 6987 6239 6993
rect 6181 6984 6193 6987
rect 5675 6956 6193 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 6181 6953 6193 6956
rect 6227 6953 6239 6987
rect 6181 6947 6239 6953
rect 6546 6944 6552 6996
rect 6604 6984 6610 6996
rect 7009 6987 7067 6993
rect 7009 6984 7021 6987
rect 6604 6956 7021 6984
rect 6604 6944 6610 6956
rect 7009 6953 7021 6956
rect 7055 6953 7067 6987
rect 7009 6947 7067 6953
rect 7558 6944 7564 6996
rect 7616 6944 7622 6996
rect 10226 6944 10232 6996
rect 10284 6944 10290 6996
rect 12342 6944 12348 6996
rect 12400 6944 12406 6996
rect 13170 6944 13176 6996
rect 13228 6984 13234 6996
rect 13357 6987 13415 6993
rect 13357 6984 13369 6987
rect 13228 6956 13369 6984
rect 13228 6944 13234 6956
rect 13357 6953 13369 6956
rect 13403 6953 13415 6987
rect 13357 6947 13415 6953
rect 5534 6876 5540 6928
rect 5592 6916 5598 6928
rect 6089 6919 6147 6925
rect 6089 6916 6101 6919
rect 5592 6888 6101 6916
rect 5592 6876 5598 6888
rect 6089 6885 6101 6888
rect 6135 6885 6147 6919
rect 6089 6879 6147 6885
rect 7190 6876 7196 6928
rect 7248 6876 7254 6928
rect 7282 6876 7288 6928
rect 7340 6916 7346 6928
rect 7377 6919 7435 6925
rect 7377 6916 7389 6919
rect 7340 6888 7389 6916
rect 7340 6876 7346 6888
rect 7377 6885 7389 6888
rect 7423 6885 7435 6919
rect 7377 6879 7435 6885
rect 9950 6876 9956 6928
rect 10008 6916 10014 6928
rect 10413 6919 10471 6925
rect 10413 6916 10425 6919
rect 10008 6888 10425 6916
rect 10008 6876 10014 6888
rect 10413 6885 10425 6888
rect 10459 6885 10471 6919
rect 10413 6879 10471 6885
rect 13538 6876 13544 6928
rect 13596 6876 13602 6928
rect 4632 6820 5488 6848
rect 4505 6811 4563 6817
rect 5810 6808 5816 6860
rect 5868 6808 5874 6860
rect 5994 6808 6000 6860
rect 6052 6808 6058 6860
rect 8386 6808 8392 6860
rect 8444 6848 8450 6860
rect 8674 6851 8732 6857
rect 8674 6848 8686 6851
rect 8444 6820 8686 6848
rect 8444 6808 8450 6820
rect 8674 6817 8686 6820
rect 8720 6817 8732 6851
rect 8674 6811 8732 6817
rect 8938 6808 8944 6860
rect 8996 6808 9002 6860
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6848 10839 6851
rect 10870 6848 10876 6860
rect 10827 6820 10876 6848
rect 10827 6817 10839 6820
rect 10781 6811 10839 6817
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 10962 6808 10968 6860
rect 11020 6808 11026 6860
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11221 6851 11279 6857
rect 11221 6848 11233 6851
rect 11112 6820 11233 6848
rect 11112 6808 11118 6820
rect 11221 6817 11233 6820
rect 11267 6817 11279 6851
rect 11221 6811 11279 6817
rect 12986 6808 12992 6860
rect 13044 6848 13050 6860
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13044 6820 13737 6848
rect 13044 6808 13050 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 13725 6811 13783 6817
rect 4246 6740 4252 6792
rect 4304 6740 4310 6792
rect 5442 6740 5448 6792
rect 5500 6780 5506 6792
rect 6365 6783 6423 6789
rect 6365 6780 6377 6783
rect 5500 6752 6377 6780
rect 5500 6740 5506 6752
rect 6365 6749 6377 6752
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 4154 6712 4160 6724
rect 4080 6684 4160 6712
rect 4154 6672 4160 6684
rect 4212 6672 4218 6724
rect 5534 6644 5540 6656
rect 3712 6616 5540 6644
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 10410 6604 10416 6656
rect 10468 6604 10474 6656
rect 552 6554 23368 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 23368 6554
rect 552 6480 23368 6502
rect 3418 6400 3424 6452
rect 3476 6400 3482 6452
rect 3789 6443 3847 6449
rect 3789 6409 3801 6443
rect 3835 6440 3847 6443
rect 4062 6440 4068 6452
rect 3835 6412 4068 6440
rect 3835 6409 3847 6412
rect 3789 6403 3847 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 5994 6440 6000 6452
rect 4387 6412 6000 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3292 6208 3433 6236
rect 3292 6196 3298 6208
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3421 6199 3479 6205
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6236 3755 6239
rect 3973 6239 4031 6245
rect 3973 6236 3985 6239
rect 3743 6208 3985 6236
rect 3743 6205 3755 6208
rect 3697 6199 3755 6205
rect 3973 6205 3985 6208
rect 4019 6236 4031 6239
rect 4154 6236 4160 6248
rect 4019 6208 4160 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 4356 6236 4384 6403
rect 5994 6400 6000 6412
rect 6052 6400 6058 6452
rect 10318 6400 10324 6452
rect 10376 6440 10382 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 10376 6412 10425 6440
rect 10376 6400 10382 6412
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 10413 6403 10471 6409
rect 5718 6264 5724 6316
rect 5776 6304 5782 6316
rect 6822 6304 6828 6316
rect 5776 6276 6828 6304
rect 5776 6264 5782 6276
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 4295 6208 4384 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 3252 6100 3280 6196
rect 3326 6128 3332 6180
rect 3384 6168 3390 6180
rect 3513 6171 3571 6177
rect 3513 6168 3525 6171
rect 3384 6140 3525 6168
rect 3384 6128 3390 6140
rect 3513 6137 3525 6140
rect 3559 6168 3571 6171
rect 4264 6168 4292 6199
rect 5074 6196 5080 6248
rect 5132 6236 5138 6248
rect 5454 6239 5512 6245
rect 5454 6236 5466 6239
rect 5132 6208 5466 6236
rect 5132 6196 5138 6208
rect 5454 6205 5466 6208
rect 5500 6205 5512 6239
rect 5454 6199 5512 6205
rect 10597 6239 10655 6245
rect 10597 6205 10609 6239
rect 10643 6236 10655 6239
rect 10686 6236 10692 6248
rect 10643 6208 10692 6236
rect 10643 6205 10655 6208
rect 10597 6199 10655 6205
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 3559 6140 4292 6168
rect 10781 6171 10839 6177
rect 3559 6137 3571 6140
rect 3513 6131 3571 6137
rect 10781 6137 10793 6171
rect 10827 6168 10839 6171
rect 11606 6168 11612 6180
rect 10827 6140 11612 6168
rect 10827 6137 10839 6140
rect 10781 6131 10839 6137
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 4157 6103 4215 6109
rect 4157 6100 4169 6103
rect 3252 6072 4169 6100
rect 4157 6069 4169 6072
rect 4203 6100 4215 6103
rect 5810 6100 5816 6112
rect 4203 6072 5816 6100
rect 4203 6069 4215 6072
rect 4157 6063 4215 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 552 6010 23368 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 23368 6010
rect 552 5936 23368 5958
rect 5261 5899 5319 5905
rect 5261 5865 5273 5899
rect 5307 5896 5319 5899
rect 5810 5896 5816 5908
rect 5307 5868 5816 5896
rect 5307 5865 5319 5868
rect 5261 5859 5319 5865
rect 5810 5856 5816 5868
rect 5868 5856 5874 5908
rect 3510 5788 3516 5840
rect 3568 5828 3574 5840
rect 4126 5831 4184 5837
rect 4126 5828 4138 5831
rect 3568 5800 4138 5828
rect 3568 5788 3574 5800
rect 4126 5797 4138 5800
rect 4172 5797 4184 5831
rect 4126 5791 4184 5797
rect 3881 5763 3939 5769
rect 3881 5729 3893 5763
rect 3927 5760 3939 5763
rect 5718 5760 5724 5772
rect 3927 5732 5724 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 552 5466 23368 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 23368 5466
rect 552 5392 23368 5414
rect 552 4922 23368 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 23368 4922
rect 552 4848 23368 4870
rect 552 4378 23368 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 23368 4378
rect 552 4304 23368 4326
rect 22738 4088 22744 4140
rect 22796 4088 22802 4140
rect 22922 3952 22928 4004
rect 22980 3952 22986 4004
rect 552 3834 23368 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 23368 3834
rect 552 3760 23368 3782
rect 552 3290 23368 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 23368 3290
rect 552 3216 23368 3238
rect 552 2746 23368 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 23368 2746
rect 552 2672 23368 2694
rect 552 2202 23368 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 23368 2202
rect 552 2128 23368 2150
rect 552 1658 23368 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 23368 1658
rect 552 1584 23368 1606
rect 552 1114 23368 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 23368 1114
rect 552 1040 23368 1062
rect 552 570 23368 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 23368 570
rect 552 496 23368 518
<< via1 >>
rect 4322 23366 4374 23418
rect 4386 23366 4438 23418
rect 4450 23366 4502 23418
rect 4514 23366 4566 23418
rect 4578 23366 4630 23418
rect 4712 23196 4764 23248
rect 1768 23171 1820 23180
rect 1768 23137 1777 23171
rect 1777 23137 1811 23171
rect 1811 23137 1820 23171
rect 1768 23128 1820 23137
rect 10508 23196 10560 23248
rect 5356 23128 5408 23180
rect 6460 23171 6512 23180
rect 6460 23137 6469 23171
rect 6469 23137 6503 23171
rect 6503 23137 6512 23171
rect 6460 23128 6512 23137
rect 6920 23128 6972 23180
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 8668 23171 8720 23180
rect 8668 23137 8677 23171
rect 8677 23137 8711 23171
rect 8711 23137 8720 23171
rect 8668 23128 8720 23137
rect 8852 23171 8904 23180
rect 8852 23137 8861 23171
rect 8861 23137 8895 23171
rect 8895 23137 8904 23171
rect 8852 23128 8904 23137
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 16488 23171 16540 23180
rect 16488 23137 16497 23171
rect 16497 23137 16531 23171
rect 16531 23137 16540 23171
rect 16488 23128 16540 23137
rect 7472 23060 7524 23112
rect 8300 23060 8352 23112
rect 9220 23060 9272 23112
rect 9496 23060 9548 23112
rect 10140 23060 10192 23112
rect 15292 23060 15344 23112
rect 18880 23239 18932 23248
rect 18880 23205 18905 23239
rect 18905 23205 18932 23239
rect 18880 23196 18932 23205
rect 20076 23196 20128 23248
rect 20260 23196 20312 23248
rect 20904 23196 20956 23248
rect 19064 23128 19116 23180
rect 19248 23128 19300 23180
rect 19432 23171 19484 23180
rect 19432 23137 19441 23171
rect 19441 23137 19475 23171
rect 19475 23137 19484 23171
rect 19432 23128 19484 23137
rect 21180 23128 21232 23180
rect 21456 23171 21508 23180
rect 21456 23137 21465 23171
rect 21465 23137 21499 23171
rect 21499 23137 21508 23171
rect 21456 23128 21508 23137
rect 22284 23128 22336 23180
rect 20812 23060 20864 23112
rect 22652 23060 22704 23112
rect 8116 22992 8168 23044
rect 9036 23035 9088 23044
rect 9036 23001 9045 23035
rect 9045 23001 9079 23035
rect 9079 23001 9088 23035
rect 9036 22992 9088 23001
rect 18144 22992 18196 23044
rect 4896 22967 4948 22976
rect 4896 22933 4905 22967
rect 4905 22933 4939 22967
rect 4939 22933 4948 22967
rect 4896 22924 4948 22933
rect 5356 22967 5408 22976
rect 5356 22933 5365 22967
rect 5365 22933 5399 22967
rect 5399 22933 5408 22967
rect 5356 22924 5408 22933
rect 11336 22967 11388 22976
rect 11336 22933 11345 22967
rect 11345 22933 11379 22967
rect 11379 22933 11388 22967
rect 11336 22924 11388 22933
rect 14924 22924 14976 22976
rect 16672 22967 16724 22976
rect 16672 22933 16681 22967
rect 16681 22933 16715 22967
rect 16715 22933 16724 22967
rect 16672 22924 16724 22933
rect 17960 22924 18012 22976
rect 20720 22992 20772 23044
rect 19064 22967 19116 22976
rect 19064 22933 19073 22967
rect 19073 22933 19107 22967
rect 19107 22933 19116 22967
rect 19064 22924 19116 22933
rect 19156 22967 19208 22976
rect 19156 22933 19165 22967
rect 19165 22933 19199 22967
rect 19199 22933 19208 22967
rect 19156 22924 19208 22933
rect 20168 22924 20220 22976
rect 21180 22924 21232 22976
rect 21640 22967 21692 22976
rect 21640 22933 21649 22967
rect 21649 22933 21683 22967
rect 21683 22933 21692 22967
rect 21640 22924 21692 22933
rect 3662 22822 3714 22874
rect 3726 22822 3778 22874
rect 3790 22822 3842 22874
rect 3854 22822 3906 22874
rect 3918 22822 3970 22874
rect 4712 22695 4764 22704
rect 4712 22661 4721 22695
rect 4721 22661 4755 22695
rect 4755 22661 4764 22695
rect 4712 22652 4764 22661
rect 4896 22652 4948 22704
rect 6920 22720 6972 22772
rect 8208 22720 8260 22772
rect 8668 22720 8720 22772
rect 9312 22720 9364 22772
rect 12164 22720 12216 22772
rect 12808 22763 12860 22772
rect 12808 22729 12817 22763
rect 12817 22729 12851 22763
rect 12851 22729 12860 22763
rect 12808 22720 12860 22729
rect 15200 22720 15252 22772
rect 8484 22652 8536 22704
rect 4804 22516 4856 22568
rect 4252 22448 4304 22500
rect 5356 22516 5408 22568
rect 5908 22559 5960 22568
rect 5908 22525 5917 22559
rect 5917 22525 5951 22559
rect 5951 22525 5960 22559
rect 5908 22516 5960 22525
rect 6368 22559 6420 22568
rect 6368 22525 6377 22559
rect 6377 22525 6411 22559
rect 6411 22525 6420 22559
rect 6368 22516 6420 22525
rect 7472 22559 7524 22568
rect 7472 22525 7481 22559
rect 7481 22525 7515 22559
rect 7515 22525 7524 22559
rect 7472 22516 7524 22525
rect 7564 22559 7616 22568
rect 7564 22525 7573 22559
rect 7573 22525 7607 22559
rect 7607 22525 7616 22559
rect 7564 22516 7616 22525
rect 8208 22584 8260 22636
rect 7196 22448 7248 22500
rect 8024 22516 8076 22568
rect 7564 22380 7616 22432
rect 8300 22448 8352 22500
rect 8576 22380 8628 22432
rect 8760 22559 8812 22568
rect 8760 22525 8769 22559
rect 8769 22525 8803 22559
rect 8803 22525 8812 22559
rect 8760 22516 8812 22525
rect 8852 22559 8904 22568
rect 8852 22525 8861 22559
rect 8861 22525 8895 22559
rect 8895 22525 8904 22559
rect 8852 22516 8904 22525
rect 9036 22652 9088 22704
rect 11980 22652 12032 22704
rect 9312 22559 9364 22568
rect 9312 22525 9321 22559
rect 9321 22525 9355 22559
rect 9355 22525 9364 22559
rect 9312 22516 9364 22525
rect 9496 22559 9548 22568
rect 9496 22525 9505 22559
rect 9505 22525 9539 22559
rect 9539 22525 9548 22559
rect 9496 22516 9548 22525
rect 9588 22559 9640 22568
rect 9588 22525 9597 22559
rect 9597 22525 9631 22559
rect 9631 22525 9640 22559
rect 9588 22516 9640 22525
rect 11704 22584 11756 22636
rect 9864 22491 9916 22500
rect 9864 22457 9873 22491
rect 9873 22457 9907 22491
rect 9907 22457 9916 22491
rect 9864 22448 9916 22457
rect 10600 22559 10652 22568
rect 10600 22525 10610 22559
rect 10610 22525 10644 22559
rect 10644 22525 10652 22559
rect 10600 22516 10652 22525
rect 12900 22652 12952 22704
rect 13636 22652 13688 22704
rect 15568 22652 15620 22704
rect 17224 22720 17276 22772
rect 21456 22720 21508 22772
rect 21548 22763 21600 22772
rect 21548 22729 21557 22763
rect 21557 22729 21591 22763
rect 21591 22729 21600 22763
rect 21548 22720 21600 22729
rect 16488 22652 16540 22704
rect 12348 22491 12400 22500
rect 12348 22457 12357 22491
rect 12357 22457 12391 22491
rect 12391 22457 12400 22491
rect 12348 22448 12400 22457
rect 13544 22559 13596 22568
rect 13544 22525 13553 22559
rect 13553 22525 13587 22559
rect 13587 22525 13596 22559
rect 13544 22516 13596 22525
rect 13636 22559 13688 22568
rect 13636 22525 13646 22559
rect 13646 22525 13680 22559
rect 13680 22525 13688 22559
rect 13636 22516 13688 22525
rect 13268 22448 13320 22500
rect 16580 22516 16632 22568
rect 17224 22584 17276 22636
rect 17960 22627 18012 22636
rect 17960 22593 17969 22627
rect 17969 22593 18003 22627
rect 18003 22593 18012 22627
rect 17960 22584 18012 22593
rect 19248 22652 19300 22704
rect 18880 22584 18932 22636
rect 19156 22627 19208 22636
rect 19156 22593 19165 22627
rect 19165 22593 19199 22627
rect 19199 22593 19208 22627
rect 19156 22584 19208 22593
rect 18144 22559 18196 22568
rect 18144 22525 18153 22559
rect 18153 22525 18187 22559
rect 18187 22525 18196 22559
rect 18144 22516 18196 22525
rect 18788 22516 18840 22568
rect 19800 22559 19852 22568
rect 19800 22525 19809 22559
rect 19809 22525 19843 22559
rect 19843 22525 19852 22559
rect 20168 22559 20220 22568
rect 19800 22516 19852 22525
rect 20168 22525 20177 22559
rect 20177 22525 20211 22559
rect 20211 22525 20220 22559
rect 20168 22516 20220 22525
rect 20260 22559 20312 22568
rect 20260 22525 20269 22559
rect 20269 22525 20303 22559
rect 20303 22525 20312 22559
rect 20260 22516 20312 22525
rect 20904 22652 20956 22704
rect 21824 22652 21876 22704
rect 20812 22627 20864 22636
rect 20812 22593 20821 22627
rect 20821 22593 20855 22627
rect 20855 22593 20864 22627
rect 20812 22584 20864 22593
rect 21364 22584 21416 22636
rect 21640 22584 21692 22636
rect 20720 22559 20772 22568
rect 20720 22525 20729 22559
rect 20729 22525 20763 22559
rect 20763 22525 20772 22559
rect 20720 22516 20772 22525
rect 21180 22559 21232 22568
rect 21180 22525 21189 22559
rect 21189 22525 21223 22559
rect 21223 22525 21232 22559
rect 21180 22516 21232 22525
rect 21272 22559 21324 22568
rect 21272 22525 21281 22559
rect 21281 22525 21315 22559
rect 21315 22525 21324 22559
rect 21272 22516 21324 22525
rect 21456 22559 21508 22568
rect 21456 22525 21465 22559
rect 21465 22525 21499 22559
rect 21499 22525 21508 22559
rect 21456 22516 21508 22525
rect 15292 22491 15344 22500
rect 15292 22457 15301 22491
rect 15301 22457 15335 22491
rect 15335 22457 15344 22491
rect 15292 22448 15344 22457
rect 16672 22448 16724 22500
rect 8944 22380 8996 22432
rect 9312 22380 9364 22432
rect 10876 22423 10928 22432
rect 10876 22389 10885 22423
rect 10885 22389 10919 22423
rect 10919 22389 10928 22423
rect 10876 22380 10928 22389
rect 11060 22423 11112 22432
rect 11060 22389 11069 22423
rect 11069 22389 11103 22423
rect 11103 22389 11112 22423
rect 11060 22380 11112 22389
rect 12532 22423 12584 22432
rect 12532 22389 12557 22423
rect 12557 22389 12584 22423
rect 12532 22380 12584 22389
rect 12716 22423 12768 22432
rect 12716 22389 12725 22423
rect 12725 22389 12759 22423
rect 12759 22389 12768 22423
rect 12716 22380 12768 22389
rect 13176 22423 13228 22432
rect 13176 22389 13185 22423
rect 13185 22389 13219 22423
rect 13219 22389 13228 22423
rect 13176 22380 13228 22389
rect 13912 22423 13964 22432
rect 13912 22389 13921 22423
rect 13921 22389 13955 22423
rect 13955 22389 13964 22423
rect 13912 22380 13964 22389
rect 14372 22423 14424 22432
rect 14372 22389 14381 22423
rect 14381 22389 14415 22423
rect 14415 22389 14424 22423
rect 14372 22380 14424 22389
rect 15936 22380 15988 22432
rect 16488 22380 16540 22432
rect 17132 22448 17184 22500
rect 17316 22448 17368 22500
rect 20352 22448 20404 22500
rect 17684 22423 17736 22432
rect 17684 22389 17709 22423
rect 17709 22389 17736 22423
rect 17684 22380 17736 22389
rect 17868 22423 17920 22432
rect 17868 22389 17877 22423
rect 17877 22389 17911 22423
rect 17911 22389 17920 22423
rect 17868 22380 17920 22389
rect 20076 22380 20128 22432
rect 22100 22380 22152 22432
rect 22192 22423 22244 22432
rect 22192 22389 22201 22423
rect 22201 22389 22235 22423
rect 22235 22389 22244 22423
rect 22192 22380 22244 22389
rect 4322 22278 4374 22330
rect 4386 22278 4438 22330
rect 4450 22278 4502 22330
rect 4514 22278 4566 22330
rect 4578 22278 4630 22330
rect 4804 22219 4856 22228
rect 4804 22185 4813 22219
rect 4813 22185 4847 22219
rect 4847 22185 4856 22219
rect 4804 22176 4856 22185
rect 8944 22176 8996 22228
rect 9588 22176 9640 22228
rect 12348 22176 12400 22228
rect 4252 22108 4304 22160
rect 5632 22108 5684 22160
rect 6460 22108 6512 22160
rect 6736 22108 6788 22160
rect 9036 22108 9088 22160
rect 6828 22083 6880 22092
rect 6828 22049 6837 22083
rect 6837 22049 6871 22083
rect 6871 22049 6880 22083
rect 6828 22040 6880 22049
rect 7196 22083 7248 22092
rect 7196 22049 7205 22083
rect 7205 22049 7239 22083
rect 7239 22049 7248 22083
rect 7196 22040 7248 22049
rect 8116 22083 8168 22092
rect 8116 22049 8125 22083
rect 8125 22049 8159 22083
rect 8159 22049 8168 22083
rect 8116 22040 8168 22049
rect 9864 22040 9916 22092
rect 11152 22040 11204 22092
rect 12900 22108 12952 22160
rect 13912 22176 13964 22228
rect 15108 22176 15160 22228
rect 15568 22176 15620 22228
rect 16120 22176 16172 22228
rect 19156 22176 19208 22228
rect 20260 22176 20312 22228
rect 21180 22176 21232 22228
rect 12532 22040 12584 22092
rect 14924 22083 14976 22092
rect 14924 22049 14933 22083
rect 14933 22049 14967 22083
rect 14967 22049 14976 22083
rect 14924 22040 14976 22049
rect 4988 21972 5040 22024
rect 4712 21904 4764 21956
rect 6920 21904 6972 21956
rect 8300 21972 8352 22024
rect 8852 21972 8904 22024
rect 7472 21904 7524 21956
rect 8116 21904 8168 21956
rect 9404 22015 9456 22024
rect 9404 21981 9413 22015
rect 9413 21981 9447 22015
rect 9447 21981 9456 22015
rect 9404 21972 9456 21981
rect 11244 22015 11296 22024
rect 11244 21981 11253 22015
rect 11253 21981 11287 22015
rect 11287 21981 11296 22015
rect 11244 21972 11296 21981
rect 12164 22015 12216 22024
rect 12164 21981 12173 22015
rect 12173 21981 12207 22015
rect 12207 21981 12216 22015
rect 12164 21972 12216 21981
rect 13544 21972 13596 22024
rect 13820 22015 13872 22024
rect 13820 21981 13829 22015
rect 13829 21981 13863 22015
rect 13863 21981 13872 22015
rect 13820 21972 13872 21981
rect 14280 21972 14332 22024
rect 15200 21972 15252 22024
rect 11060 21904 11112 21956
rect 16488 22108 16540 22160
rect 15752 22083 15804 22092
rect 15752 22049 15761 22083
rect 15761 22049 15795 22083
rect 15795 22049 15804 22083
rect 15752 22040 15804 22049
rect 16120 22083 16172 22092
rect 16120 22049 16129 22083
rect 16129 22049 16163 22083
rect 16163 22049 16172 22083
rect 16120 22040 16172 22049
rect 16212 22040 16264 22092
rect 17592 22108 17644 22160
rect 19340 22108 19392 22160
rect 20352 22108 20404 22160
rect 15660 22015 15712 22024
rect 15660 21981 15669 22015
rect 15669 21981 15703 22015
rect 15703 21981 15712 22015
rect 15660 21972 15712 21981
rect 17040 22083 17092 22092
rect 17040 22049 17049 22083
rect 17049 22049 17083 22083
rect 17083 22049 17092 22083
rect 17040 22040 17092 22049
rect 17776 22040 17828 22092
rect 17500 21972 17552 22024
rect 19064 22040 19116 22092
rect 19248 22083 19300 22092
rect 19248 22049 19257 22083
rect 19257 22049 19291 22083
rect 19291 22049 19300 22083
rect 19248 22040 19300 22049
rect 19340 21972 19392 22024
rect 20168 22083 20220 22092
rect 20168 22049 20177 22083
rect 20177 22049 20211 22083
rect 20211 22049 20220 22083
rect 20168 22040 20220 22049
rect 20812 22108 20864 22160
rect 21364 22108 21416 22160
rect 21456 22040 21508 22092
rect 22100 22176 22152 22228
rect 22652 22151 22704 22160
rect 22652 22117 22661 22151
rect 22661 22117 22695 22151
rect 22695 22117 22704 22151
rect 22652 22108 22704 22117
rect 21732 22015 21784 22024
rect 21732 21981 21741 22015
rect 21741 21981 21775 22015
rect 21775 21981 21784 22015
rect 21732 21972 21784 21981
rect 22192 22083 22244 22092
rect 22192 22049 22201 22083
rect 22201 22049 22235 22083
rect 22235 22049 22244 22083
rect 22192 22040 22244 22049
rect 22376 22083 22428 22092
rect 22376 22049 22385 22083
rect 22385 22049 22419 22083
rect 22419 22049 22428 22083
rect 22376 22040 22428 22049
rect 19708 21904 19760 21956
rect 21640 21904 21692 21956
rect 22284 22015 22336 22024
rect 22284 21981 22293 22015
rect 22293 21981 22327 22015
rect 22327 21981 22336 22015
rect 22284 21972 22336 21981
rect 5448 21836 5500 21888
rect 8852 21836 8904 21888
rect 9312 21836 9364 21888
rect 13912 21879 13964 21888
rect 13912 21845 13921 21879
rect 13921 21845 13955 21879
rect 13955 21845 13964 21879
rect 13912 21836 13964 21845
rect 14188 21836 14240 21888
rect 17408 21836 17460 21888
rect 17684 21836 17736 21888
rect 18696 21879 18748 21888
rect 18696 21845 18705 21879
rect 18705 21845 18739 21879
rect 18739 21845 18748 21879
rect 18696 21836 18748 21845
rect 18788 21836 18840 21888
rect 20536 21879 20588 21888
rect 20536 21845 20545 21879
rect 20545 21845 20579 21879
rect 20579 21845 20588 21879
rect 20536 21836 20588 21845
rect 20996 21836 21048 21888
rect 3662 21734 3714 21786
rect 3726 21734 3778 21786
rect 3790 21734 3842 21786
rect 3854 21734 3906 21786
rect 3918 21734 3970 21786
rect 5448 21632 5500 21684
rect 6828 21564 6880 21616
rect 7656 21632 7708 21684
rect 8760 21632 8812 21684
rect 12808 21632 12860 21684
rect 15108 21632 15160 21684
rect 6276 21428 6328 21480
rect 6736 21471 6788 21480
rect 6736 21437 6745 21471
rect 6745 21437 6779 21471
rect 6779 21437 6788 21471
rect 6736 21428 6788 21437
rect 6828 21428 6880 21480
rect 7380 21360 7432 21412
rect 4712 21292 4764 21344
rect 6828 21292 6880 21344
rect 7656 21471 7708 21480
rect 7656 21437 7665 21471
rect 7665 21437 7699 21471
rect 7699 21437 7708 21471
rect 7656 21428 7708 21437
rect 8208 21564 8260 21616
rect 8024 21471 8076 21480
rect 8024 21437 8033 21471
rect 8033 21437 8067 21471
rect 8067 21437 8076 21471
rect 8024 21428 8076 21437
rect 8300 21428 8352 21480
rect 8576 21428 8628 21480
rect 8668 21471 8720 21480
rect 8668 21437 8677 21471
rect 8677 21437 8711 21471
rect 8711 21437 8720 21471
rect 8668 21428 8720 21437
rect 8944 21471 8996 21480
rect 8944 21437 8953 21471
rect 8953 21437 8987 21471
rect 8987 21437 8996 21471
rect 8944 21428 8996 21437
rect 9220 21471 9272 21480
rect 9220 21437 9229 21471
rect 9229 21437 9263 21471
rect 9263 21437 9272 21471
rect 9220 21428 9272 21437
rect 10600 21496 10652 21548
rect 10876 21539 10928 21548
rect 10876 21505 10885 21539
rect 10885 21505 10919 21539
rect 10919 21505 10928 21539
rect 10876 21496 10928 21505
rect 9496 21428 9548 21480
rect 10140 21471 10192 21480
rect 10140 21437 10149 21471
rect 10149 21437 10183 21471
rect 10183 21437 10192 21471
rect 10140 21428 10192 21437
rect 10324 21471 10376 21480
rect 10324 21437 10333 21471
rect 10333 21437 10367 21471
rect 10367 21437 10376 21471
rect 10324 21428 10376 21437
rect 10416 21428 10468 21480
rect 10692 21471 10744 21480
rect 10692 21437 10701 21471
rect 10701 21437 10735 21471
rect 10735 21437 10744 21471
rect 10692 21428 10744 21437
rect 11060 21428 11112 21480
rect 11152 21428 11204 21480
rect 11704 21471 11756 21480
rect 11704 21437 11713 21471
rect 11713 21437 11747 21471
rect 11747 21437 11756 21471
rect 11704 21428 11756 21437
rect 12348 21539 12400 21548
rect 12348 21505 12357 21539
rect 12357 21505 12391 21539
rect 12391 21505 12400 21539
rect 12348 21496 12400 21505
rect 13268 21496 13320 21548
rect 14372 21539 14424 21548
rect 14372 21505 14381 21539
rect 14381 21505 14415 21539
rect 14415 21505 14424 21539
rect 14372 21496 14424 21505
rect 15016 21539 15068 21548
rect 15016 21505 15025 21539
rect 15025 21505 15059 21539
rect 15059 21505 15068 21539
rect 15016 21496 15068 21505
rect 15660 21496 15712 21548
rect 10324 21292 10376 21344
rect 11244 21360 11296 21412
rect 12164 21428 12216 21480
rect 12256 21471 12308 21480
rect 12256 21437 12265 21471
rect 12265 21437 12299 21471
rect 12299 21437 12308 21471
rect 12256 21428 12308 21437
rect 12440 21428 12492 21480
rect 12716 21428 12768 21480
rect 14188 21471 14240 21480
rect 14188 21437 14197 21471
rect 14197 21437 14231 21471
rect 14231 21437 14240 21471
rect 14188 21428 14240 21437
rect 14924 21471 14976 21480
rect 14924 21437 14933 21471
rect 14933 21437 14967 21471
rect 14967 21437 14976 21471
rect 14924 21428 14976 21437
rect 15108 21471 15160 21480
rect 15108 21437 15117 21471
rect 15117 21437 15151 21471
rect 15151 21437 15160 21471
rect 15108 21428 15160 21437
rect 13728 21360 13780 21412
rect 11152 21292 11204 21344
rect 11428 21292 11480 21344
rect 11980 21292 12032 21344
rect 13176 21292 13228 21344
rect 13360 21335 13412 21344
rect 13360 21301 13369 21335
rect 13369 21301 13403 21335
rect 13403 21301 13412 21335
rect 13360 21292 13412 21301
rect 13452 21292 13504 21344
rect 13636 21292 13688 21344
rect 17316 21632 17368 21684
rect 17408 21632 17460 21684
rect 17132 21564 17184 21616
rect 17500 21607 17552 21616
rect 17500 21573 17509 21607
rect 17509 21573 17543 21607
rect 17543 21573 17552 21607
rect 17500 21564 17552 21573
rect 17776 21496 17828 21548
rect 15384 21403 15436 21412
rect 15384 21369 15393 21403
rect 15393 21369 15427 21403
rect 15427 21369 15436 21403
rect 15384 21360 15436 21369
rect 15568 21403 15620 21412
rect 15568 21369 15577 21403
rect 15577 21369 15611 21403
rect 15611 21369 15620 21403
rect 15568 21360 15620 21369
rect 16672 21428 16724 21480
rect 17224 21471 17276 21480
rect 17224 21437 17233 21471
rect 17233 21437 17267 21471
rect 17267 21437 17276 21471
rect 17224 21428 17276 21437
rect 17316 21471 17368 21480
rect 17316 21437 17325 21471
rect 17325 21437 17359 21471
rect 17359 21437 17368 21471
rect 17316 21428 17368 21437
rect 17684 21428 17736 21480
rect 18696 21632 18748 21684
rect 21732 21632 21784 21684
rect 18052 21539 18104 21548
rect 18052 21505 18061 21539
rect 18061 21505 18095 21539
rect 18095 21505 18104 21539
rect 18052 21496 18104 21505
rect 17040 21360 17092 21412
rect 16764 21335 16816 21344
rect 16764 21301 16773 21335
rect 16773 21301 16807 21335
rect 16807 21301 16816 21335
rect 16764 21292 16816 21301
rect 18236 21403 18288 21412
rect 18236 21369 18245 21403
rect 18245 21369 18279 21403
rect 18279 21369 18288 21403
rect 18236 21360 18288 21369
rect 21548 21564 21600 21616
rect 22284 21496 22336 21548
rect 20996 21471 21048 21480
rect 20996 21437 21005 21471
rect 21005 21437 21039 21471
rect 21039 21437 21048 21471
rect 20996 21428 21048 21437
rect 21272 21428 21324 21480
rect 20076 21335 20128 21344
rect 20076 21301 20085 21335
rect 20085 21301 20119 21335
rect 20119 21301 20128 21335
rect 20076 21292 20128 21301
rect 20996 21292 21048 21344
rect 21272 21335 21324 21344
rect 21272 21301 21281 21335
rect 21281 21301 21315 21335
rect 21315 21301 21324 21335
rect 21272 21292 21324 21301
rect 4322 21190 4374 21242
rect 4386 21190 4438 21242
rect 4450 21190 4502 21242
rect 4514 21190 4566 21242
rect 4578 21190 4630 21242
rect 6736 21088 6788 21140
rect 8024 21088 8076 21140
rect 5908 21020 5960 21072
rect 4712 20952 4764 21004
rect 5632 20995 5684 21004
rect 5632 20961 5641 20995
rect 5641 20961 5675 20995
rect 5675 20961 5684 20995
rect 5632 20952 5684 20961
rect 6368 20884 6420 20936
rect 7012 20927 7064 20936
rect 7012 20893 7021 20927
rect 7021 20893 7055 20927
rect 7055 20893 7064 20927
rect 7012 20884 7064 20893
rect 7380 20995 7432 21004
rect 7380 20961 7389 20995
rect 7389 20961 7423 20995
rect 7423 20961 7432 20995
rect 7380 20952 7432 20961
rect 8300 20952 8352 21004
rect 9220 21020 9272 21072
rect 9588 21088 9640 21140
rect 8576 20952 8628 21004
rect 9772 21020 9824 21072
rect 8116 20884 8168 20936
rect 6736 20816 6788 20868
rect 8760 20816 8812 20868
rect 9220 20884 9272 20936
rect 9680 20995 9732 21004
rect 9680 20961 9689 20995
rect 9689 20961 9723 20995
rect 9723 20961 9732 20995
rect 9680 20952 9732 20961
rect 10416 21131 10468 21140
rect 10416 21097 10425 21131
rect 10425 21097 10459 21131
rect 10459 21097 10468 21131
rect 10416 21088 10468 21097
rect 13636 21088 13688 21140
rect 10232 20995 10284 21004
rect 10232 20961 10241 20995
rect 10241 20961 10275 20995
rect 10275 20961 10284 20995
rect 10232 20952 10284 20961
rect 10508 20995 10560 21004
rect 10508 20961 10517 20995
rect 10517 20961 10551 20995
rect 10551 20961 10560 20995
rect 10508 20952 10560 20961
rect 10416 20884 10468 20936
rect 9404 20816 9456 20868
rect 13728 20952 13780 21004
rect 13820 20952 13872 21004
rect 15292 21088 15344 21140
rect 16672 21131 16724 21140
rect 16672 21097 16681 21131
rect 16681 21097 16715 21131
rect 16715 21097 16724 21131
rect 16672 21088 16724 21097
rect 17868 21088 17920 21140
rect 18052 21131 18104 21140
rect 18052 21097 18061 21131
rect 18061 21097 18095 21131
rect 18095 21097 18104 21131
rect 18052 21088 18104 21097
rect 15016 21020 15068 21072
rect 15200 20952 15252 21004
rect 15936 20995 15988 21004
rect 15936 20961 15945 20995
rect 15945 20961 15979 20995
rect 15979 20961 15988 20995
rect 15936 20952 15988 20961
rect 21272 21088 21324 21140
rect 13636 20884 13688 20936
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 15384 20884 15436 20936
rect 16580 20952 16632 21004
rect 17132 20952 17184 21004
rect 17500 20952 17552 21004
rect 18236 20952 18288 21004
rect 20076 20995 20128 21004
rect 20076 20961 20085 20995
rect 20085 20961 20119 20995
rect 20119 20961 20128 20995
rect 20076 20952 20128 20961
rect 17316 20884 17368 20936
rect 20352 20995 20404 21004
rect 20352 20961 20361 20995
rect 20361 20961 20395 20995
rect 20395 20961 20404 20995
rect 20352 20952 20404 20961
rect 20996 21020 21048 21072
rect 21548 21020 21600 21072
rect 22284 20952 22336 21004
rect 6092 20748 6144 20800
rect 6368 20791 6420 20800
rect 6368 20757 6377 20791
rect 6377 20757 6411 20791
rect 6411 20757 6420 20791
rect 6368 20748 6420 20757
rect 6644 20748 6696 20800
rect 7840 20791 7892 20800
rect 7840 20757 7849 20791
rect 7849 20757 7883 20791
rect 7883 20757 7892 20791
rect 7840 20748 7892 20757
rect 8300 20748 8352 20800
rect 9220 20748 9272 20800
rect 9588 20791 9640 20800
rect 9588 20757 9597 20791
rect 9597 20757 9631 20791
rect 9631 20757 9640 20791
rect 9588 20748 9640 20757
rect 10692 20748 10744 20800
rect 12624 20748 12676 20800
rect 16212 20816 16264 20868
rect 20352 20816 20404 20868
rect 18696 20748 18748 20800
rect 19524 20748 19576 20800
rect 20628 20791 20680 20800
rect 20628 20757 20637 20791
rect 20637 20757 20671 20791
rect 20671 20757 20680 20791
rect 20628 20748 20680 20757
rect 20720 20791 20772 20800
rect 20720 20757 20729 20791
rect 20729 20757 20763 20791
rect 20763 20757 20772 20791
rect 20720 20748 20772 20757
rect 21272 20791 21324 20800
rect 21272 20757 21281 20791
rect 21281 20757 21315 20791
rect 21315 20757 21324 20791
rect 21272 20748 21324 20757
rect 3662 20646 3714 20698
rect 3726 20646 3778 20698
rect 3790 20646 3842 20698
rect 3854 20646 3906 20698
rect 3918 20646 3970 20698
rect 7012 20544 7064 20596
rect 20628 20587 20680 20596
rect 20628 20553 20637 20587
rect 20637 20553 20671 20587
rect 20671 20553 20680 20587
rect 20628 20544 20680 20553
rect 7656 20476 7708 20528
rect 11612 20476 11664 20528
rect 4252 20340 4304 20392
rect 4620 20383 4672 20392
rect 4620 20349 4629 20383
rect 4629 20349 4663 20383
rect 4663 20349 4672 20383
rect 4620 20340 4672 20349
rect 4804 20383 4856 20392
rect 4804 20349 4813 20383
rect 4813 20349 4847 20383
rect 4847 20349 4856 20383
rect 4804 20340 4856 20349
rect 5080 20340 5132 20392
rect 9680 20408 9732 20460
rect 5632 20383 5684 20392
rect 5632 20349 5641 20383
rect 5641 20349 5675 20383
rect 5675 20349 5684 20383
rect 5632 20340 5684 20349
rect 6092 20383 6144 20392
rect 6092 20349 6101 20383
rect 6101 20349 6135 20383
rect 6135 20349 6144 20383
rect 6092 20340 6144 20349
rect 6736 20383 6788 20392
rect 6736 20349 6745 20383
rect 6745 20349 6779 20383
rect 6779 20349 6788 20383
rect 6736 20340 6788 20349
rect 10968 20340 11020 20392
rect 11980 20383 12032 20392
rect 11980 20349 11989 20383
rect 11989 20349 12023 20383
rect 12023 20349 12032 20383
rect 11980 20340 12032 20349
rect 12624 20383 12676 20392
rect 12624 20349 12633 20383
rect 12633 20349 12667 20383
rect 12667 20349 12676 20383
rect 12624 20340 12676 20349
rect 13084 20340 13136 20392
rect 19064 20340 19116 20392
rect 19524 20383 19576 20392
rect 19524 20349 19533 20383
rect 19533 20349 19567 20383
rect 19567 20349 19576 20383
rect 19524 20340 19576 20349
rect 20720 20408 20772 20460
rect 21272 20408 21324 20460
rect 20628 20383 20680 20392
rect 20628 20349 20637 20383
rect 20637 20349 20671 20383
rect 20671 20349 20680 20383
rect 20628 20340 20680 20349
rect 20812 20340 20864 20392
rect 21456 20383 21508 20392
rect 21456 20349 21465 20383
rect 21465 20349 21499 20383
rect 21499 20349 21508 20383
rect 21456 20340 21508 20349
rect 22652 20340 22704 20392
rect 5172 20272 5224 20324
rect 18972 20272 19024 20324
rect 21824 20315 21876 20324
rect 21824 20281 21833 20315
rect 21833 20281 21867 20315
rect 21867 20281 21876 20315
rect 21824 20272 21876 20281
rect 22468 20315 22520 20324
rect 22468 20281 22477 20315
rect 22477 20281 22511 20315
rect 22511 20281 22520 20315
rect 22468 20272 22520 20281
rect 4252 20247 4304 20256
rect 4252 20213 4261 20247
rect 4261 20213 4295 20247
rect 4295 20213 4304 20247
rect 4252 20204 4304 20213
rect 6000 20247 6052 20256
rect 6000 20213 6009 20247
rect 6009 20213 6043 20247
rect 6043 20213 6052 20247
rect 6000 20204 6052 20213
rect 12532 20204 12584 20256
rect 12992 20204 13044 20256
rect 19708 20204 19760 20256
rect 20904 20247 20956 20256
rect 20904 20213 20913 20247
rect 20913 20213 20947 20247
rect 20947 20213 20956 20247
rect 20904 20204 20956 20213
rect 21916 20247 21968 20256
rect 21916 20213 21925 20247
rect 21925 20213 21959 20247
rect 21959 20213 21968 20247
rect 21916 20204 21968 20213
rect 22008 20204 22060 20256
rect 4322 20102 4374 20154
rect 4386 20102 4438 20154
rect 4450 20102 4502 20154
rect 4514 20102 4566 20154
rect 4578 20102 4630 20154
rect 5080 20043 5132 20052
rect 5080 20009 5089 20043
rect 5089 20009 5123 20043
rect 5123 20009 5132 20043
rect 5080 20000 5132 20009
rect 4160 19932 4212 19984
rect 4896 19932 4948 19984
rect 5172 19907 5224 19916
rect 5172 19873 5181 19907
rect 5181 19873 5215 19907
rect 5215 19873 5224 19907
rect 5172 19864 5224 19873
rect 6000 19907 6052 19916
rect 6000 19873 6009 19907
rect 6009 19873 6043 19907
rect 6043 19873 6052 19907
rect 6000 19864 6052 19873
rect 7012 19907 7064 19916
rect 7012 19873 7021 19907
rect 7021 19873 7055 19907
rect 7055 19873 7064 19907
rect 7012 19864 7064 19873
rect 10508 19864 10560 19916
rect 10968 19932 11020 19984
rect 15936 20000 15988 20052
rect 12348 19932 12400 19984
rect 14556 19932 14608 19984
rect 17960 20000 18012 20052
rect 18236 20000 18288 20052
rect 21456 20043 21508 20052
rect 21456 20009 21465 20043
rect 21465 20009 21499 20043
rect 21499 20009 21508 20043
rect 21456 20000 21508 20009
rect 11152 19864 11204 19916
rect 12072 19864 12124 19916
rect 12256 19864 12308 19916
rect 12624 19864 12676 19916
rect 6092 19839 6144 19848
rect 6092 19805 6101 19839
rect 6101 19805 6135 19839
rect 6135 19805 6144 19839
rect 6092 19796 6144 19805
rect 7564 19796 7616 19848
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 13084 19796 13136 19805
rect 13912 19864 13964 19916
rect 16764 19864 16816 19916
rect 17776 19975 17828 19984
rect 17776 19941 17801 19975
rect 17801 19941 17828 19975
rect 17776 19932 17828 19941
rect 18144 19932 18196 19984
rect 18512 19932 18564 19984
rect 19064 19975 19116 19984
rect 19064 19941 19073 19975
rect 19073 19941 19107 19975
rect 19107 19941 19116 19975
rect 19064 19932 19116 19941
rect 4344 19771 4396 19780
rect 4344 19737 4353 19771
rect 4353 19737 4387 19771
rect 4387 19737 4396 19771
rect 4344 19728 4396 19737
rect 4252 19660 4304 19712
rect 7104 19728 7156 19780
rect 4804 19660 4856 19712
rect 5540 19703 5592 19712
rect 5540 19669 5549 19703
rect 5549 19669 5583 19703
rect 5583 19669 5592 19703
rect 5540 19660 5592 19669
rect 13544 19771 13596 19780
rect 13544 19737 13553 19771
rect 13553 19737 13587 19771
rect 13587 19737 13596 19771
rect 13544 19728 13596 19737
rect 16856 19771 16908 19780
rect 16856 19737 16865 19771
rect 16865 19737 16899 19771
rect 16899 19737 16908 19771
rect 16856 19728 16908 19737
rect 18972 19907 19024 19916
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 18972 19873 18981 19907
rect 18981 19873 19015 19907
rect 19015 19873 19024 19907
rect 18972 19864 19024 19873
rect 19524 19864 19576 19916
rect 19708 19907 19760 19916
rect 19708 19873 19717 19907
rect 19717 19873 19751 19907
rect 19751 19873 19760 19907
rect 19708 19864 19760 19873
rect 20352 19932 20404 19984
rect 21180 19932 21232 19984
rect 22008 19932 22060 19984
rect 20168 19907 20220 19916
rect 20168 19873 20177 19907
rect 20177 19873 20211 19907
rect 20211 19873 20220 19907
rect 20168 19864 20220 19873
rect 20536 19907 20588 19916
rect 20536 19873 20545 19907
rect 20545 19873 20579 19907
rect 20579 19873 20588 19907
rect 20536 19864 20588 19873
rect 20720 19864 20772 19916
rect 18696 19728 18748 19780
rect 19984 19839 20036 19848
rect 19984 19805 19993 19839
rect 19993 19805 20027 19839
rect 20027 19805 20036 19839
rect 19984 19796 20036 19805
rect 21272 19796 21324 19848
rect 21916 19839 21968 19848
rect 21916 19805 21925 19839
rect 21925 19805 21959 19839
rect 21959 19805 21968 19839
rect 21916 19796 21968 19805
rect 22376 19907 22428 19916
rect 22376 19873 22385 19907
rect 22385 19873 22419 19907
rect 22419 19873 22428 19907
rect 22376 19864 22428 19873
rect 22744 19864 22796 19916
rect 22836 19796 22888 19848
rect 23020 19839 23072 19848
rect 23020 19805 23029 19839
rect 23029 19805 23063 19839
rect 23063 19805 23072 19839
rect 23020 19796 23072 19805
rect 13820 19703 13872 19712
rect 13820 19669 13829 19703
rect 13829 19669 13863 19703
rect 13863 19669 13872 19703
rect 13820 19660 13872 19669
rect 17868 19660 17920 19712
rect 18236 19660 18288 19712
rect 19524 19703 19576 19712
rect 19524 19669 19533 19703
rect 19533 19669 19567 19703
rect 19567 19669 19576 19703
rect 19524 19660 19576 19669
rect 20720 19660 20772 19712
rect 21088 19660 21140 19712
rect 22192 19660 22244 19712
rect 3662 19558 3714 19610
rect 3726 19558 3778 19610
rect 3790 19558 3842 19610
rect 3854 19558 3906 19610
rect 3918 19558 3970 19610
rect 4804 19456 4856 19508
rect 5172 19456 5224 19508
rect 9864 19456 9916 19508
rect 13084 19456 13136 19508
rect 14740 19456 14792 19508
rect 18696 19499 18748 19508
rect 18696 19465 18705 19499
rect 18705 19465 18739 19499
rect 18739 19465 18748 19499
rect 18696 19456 18748 19465
rect 22192 19499 22244 19508
rect 22192 19465 22201 19499
rect 22201 19465 22235 19499
rect 22235 19465 22244 19499
rect 22192 19456 22244 19465
rect 4160 19363 4212 19372
rect 4160 19329 4169 19363
rect 4169 19329 4203 19363
rect 4203 19329 4212 19363
rect 4160 19320 4212 19329
rect 4712 19363 4764 19372
rect 4712 19329 4721 19363
rect 4721 19329 4755 19363
rect 4755 19329 4764 19363
rect 4712 19320 4764 19329
rect 5172 19363 5224 19372
rect 5172 19329 5181 19363
rect 5181 19329 5215 19363
rect 5215 19329 5224 19363
rect 5172 19320 5224 19329
rect 7104 19363 7156 19372
rect 7104 19329 7113 19363
rect 7113 19329 7147 19363
rect 7147 19329 7156 19363
rect 7104 19320 7156 19329
rect 4252 19295 4304 19304
rect 4252 19261 4261 19295
rect 4261 19261 4295 19295
rect 4295 19261 4304 19295
rect 4252 19252 4304 19261
rect 4344 19295 4396 19304
rect 4344 19261 4353 19295
rect 4353 19261 4387 19295
rect 4387 19261 4396 19295
rect 4344 19252 4396 19261
rect 4804 19295 4856 19304
rect 4804 19261 4813 19295
rect 4813 19261 4847 19295
rect 4847 19261 4856 19295
rect 4804 19252 4856 19261
rect 5448 19252 5500 19304
rect 6000 19252 6052 19304
rect 7012 19252 7064 19304
rect 7196 19295 7248 19304
rect 7196 19261 7205 19295
rect 7205 19261 7239 19295
rect 7239 19261 7248 19295
rect 7196 19252 7248 19261
rect 7472 19252 7524 19304
rect 7840 19295 7892 19304
rect 7840 19261 7849 19295
rect 7849 19261 7883 19295
rect 7883 19261 7892 19295
rect 7840 19252 7892 19261
rect 8024 19295 8076 19304
rect 8024 19261 8033 19295
rect 8033 19261 8067 19295
rect 8067 19261 8076 19295
rect 8024 19252 8076 19261
rect 11980 19320 12032 19372
rect 12164 19431 12216 19440
rect 12164 19397 12173 19431
rect 12173 19397 12207 19431
rect 12207 19397 12216 19431
rect 12164 19388 12216 19397
rect 12992 19431 13044 19440
rect 12992 19397 13001 19431
rect 13001 19397 13035 19431
rect 13035 19397 13044 19431
rect 12992 19388 13044 19397
rect 12348 19320 12400 19372
rect 12532 19363 12584 19372
rect 12532 19329 12541 19363
rect 12541 19329 12575 19363
rect 12575 19329 12584 19363
rect 12532 19320 12584 19329
rect 13084 19320 13136 19372
rect 13912 19320 13964 19372
rect 14004 19320 14056 19372
rect 4988 19184 5040 19236
rect 6092 19227 6144 19236
rect 6092 19193 6101 19227
rect 6101 19193 6135 19227
rect 6135 19193 6144 19227
rect 6092 19184 6144 19193
rect 7932 19227 7984 19236
rect 7932 19193 7941 19227
rect 7941 19193 7975 19227
rect 7975 19193 7984 19227
rect 7932 19184 7984 19193
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 9680 19252 9732 19304
rect 10232 19295 10284 19304
rect 10232 19261 10241 19295
rect 10241 19261 10275 19295
rect 10275 19261 10284 19295
rect 10232 19252 10284 19261
rect 10876 19252 10928 19304
rect 10968 19295 11020 19304
rect 10968 19261 10977 19295
rect 10977 19261 11011 19295
rect 11011 19261 11020 19295
rect 10968 19252 11020 19261
rect 11612 19295 11664 19304
rect 11612 19261 11621 19295
rect 11621 19261 11655 19295
rect 11655 19261 11664 19295
rect 11612 19252 11664 19261
rect 12072 19295 12124 19304
rect 12072 19261 12081 19295
rect 12081 19261 12115 19295
rect 12115 19261 12124 19295
rect 12072 19252 12124 19261
rect 12256 19295 12308 19304
rect 12256 19261 12265 19295
rect 12265 19261 12299 19295
rect 12299 19261 12308 19295
rect 12256 19252 12308 19261
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 11704 19184 11756 19236
rect 13544 19252 13596 19304
rect 14188 19295 14240 19304
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 14648 19295 14700 19304
rect 14648 19261 14657 19295
rect 14657 19261 14691 19295
rect 14691 19261 14700 19295
rect 14648 19252 14700 19261
rect 14924 19295 14976 19304
rect 14924 19261 14933 19295
rect 14933 19261 14967 19295
rect 14967 19261 14976 19295
rect 14924 19252 14976 19261
rect 16856 19363 16908 19372
rect 16856 19329 16865 19363
rect 16865 19329 16899 19363
rect 16899 19329 16908 19363
rect 16856 19320 16908 19329
rect 15200 19252 15252 19304
rect 16764 19295 16816 19304
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 13820 19184 13872 19236
rect 17868 19295 17920 19304
rect 17868 19261 17877 19295
rect 17877 19261 17911 19295
rect 17911 19261 17920 19295
rect 17868 19252 17920 19261
rect 17960 19295 18012 19304
rect 17960 19261 17969 19295
rect 17969 19261 18003 19295
rect 18003 19261 18012 19295
rect 17960 19252 18012 19261
rect 18144 19295 18196 19304
rect 18144 19261 18153 19295
rect 18153 19261 18187 19295
rect 18187 19261 18196 19295
rect 18144 19252 18196 19261
rect 18236 19295 18288 19304
rect 18236 19261 18245 19295
rect 18245 19261 18279 19295
rect 18279 19261 18288 19295
rect 18236 19252 18288 19261
rect 18880 19295 18932 19304
rect 18880 19261 18889 19295
rect 18889 19261 18923 19295
rect 18923 19261 18932 19295
rect 18880 19252 18932 19261
rect 19156 19295 19208 19304
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 21088 19295 21140 19304
rect 21088 19261 21122 19295
rect 21122 19261 21140 19295
rect 19524 19184 19576 19236
rect 21088 19252 21140 19261
rect 21180 19184 21232 19236
rect 4804 19116 4856 19168
rect 5908 19116 5960 19168
rect 10324 19116 10376 19168
rect 14188 19116 14240 19168
rect 15016 19116 15068 19168
rect 17132 19159 17184 19168
rect 17132 19125 17141 19159
rect 17141 19125 17175 19159
rect 17175 19125 17184 19159
rect 17132 19116 17184 19125
rect 17960 19116 18012 19168
rect 20352 19116 20404 19168
rect 20628 19116 20680 19168
rect 22652 19295 22704 19304
rect 22652 19261 22661 19295
rect 22661 19261 22695 19295
rect 22695 19261 22704 19295
rect 22652 19252 22704 19261
rect 22836 19295 22888 19304
rect 22836 19261 22845 19295
rect 22845 19261 22879 19295
rect 22879 19261 22888 19295
rect 22836 19252 22888 19261
rect 22560 19227 22612 19236
rect 22560 19193 22569 19227
rect 22569 19193 22603 19227
rect 22603 19193 22612 19227
rect 22560 19184 22612 19193
rect 22284 19159 22336 19168
rect 22284 19125 22293 19159
rect 22293 19125 22327 19159
rect 22327 19125 22336 19159
rect 22284 19116 22336 19125
rect 4322 19014 4374 19066
rect 4386 19014 4438 19066
rect 4450 19014 4502 19066
rect 4514 19014 4566 19066
rect 4578 19014 4630 19066
rect 7472 18955 7524 18964
rect 7472 18921 7481 18955
rect 7481 18921 7515 18955
rect 7515 18921 7524 18955
rect 7472 18912 7524 18921
rect 7932 18955 7984 18964
rect 7932 18921 7941 18955
rect 7941 18921 7975 18955
rect 7975 18921 7984 18955
rect 7932 18912 7984 18921
rect 8024 18912 8076 18964
rect 5632 18844 5684 18896
rect 6828 18844 6880 18896
rect 8760 18844 8812 18896
rect 5172 18819 5224 18828
rect 5172 18785 5181 18819
rect 5181 18785 5215 18819
rect 5215 18785 5224 18819
rect 5172 18776 5224 18785
rect 5448 18819 5500 18828
rect 5448 18785 5457 18819
rect 5457 18785 5491 18819
rect 5491 18785 5500 18819
rect 5448 18776 5500 18785
rect 5816 18776 5868 18828
rect 6092 18640 6144 18692
rect 6552 18751 6604 18760
rect 6552 18717 6561 18751
rect 6561 18717 6595 18751
rect 6595 18717 6604 18751
rect 6552 18708 6604 18717
rect 6828 18708 6880 18760
rect 8484 18819 8536 18828
rect 8484 18785 8493 18819
rect 8493 18785 8527 18819
rect 8527 18785 8536 18819
rect 8484 18776 8536 18785
rect 9588 18887 9640 18896
rect 9588 18853 9597 18887
rect 9597 18853 9631 18887
rect 9631 18853 9640 18887
rect 9588 18844 9640 18853
rect 12808 18912 12860 18964
rect 14648 18912 14700 18964
rect 17684 18912 17736 18964
rect 18880 18912 18932 18964
rect 19984 18955 20036 18964
rect 19984 18921 19993 18955
rect 19993 18921 20027 18955
rect 20027 18921 20036 18955
rect 19984 18912 20036 18921
rect 21824 18912 21876 18964
rect 22560 18912 22612 18964
rect 9036 18776 9088 18828
rect 10968 18844 11020 18896
rect 6920 18640 6972 18692
rect 8116 18683 8168 18692
rect 8116 18649 8125 18683
rect 8125 18649 8159 18683
rect 8159 18649 8168 18683
rect 8116 18640 8168 18649
rect 10416 18819 10468 18828
rect 10416 18785 10425 18819
rect 10425 18785 10459 18819
rect 10459 18785 10468 18819
rect 10416 18776 10468 18785
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 7196 18572 7248 18624
rect 9864 18640 9916 18692
rect 9956 18683 10008 18692
rect 9956 18649 9965 18683
rect 9965 18649 9999 18683
rect 9999 18649 10008 18683
rect 11520 18776 11572 18828
rect 12164 18776 12216 18828
rect 13084 18819 13136 18828
rect 13084 18785 13093 18819
rect 13093 18785 13127 18819
rect 13127 18785 13136 18819
rect 13084 18776 13136 18785
rect 10876 18708 10928 18760
rect 9956 18640 10008 18649
rect 11980 18708 12032 18760
rect 12992 18708 13044 18760
rect 11796 18683 11848 18692
rect 11796 18649 11805 18683
rect 11805 18649 11839 18683
rect 11839 18649 11848 18683
rect 13820 18776 13872 18828
rect 14280 18819 14332 18828
rect 14280 18785 14289 18819
rect 14289 18785 14323 18819
rect 14323 18785 14332 18819
rect 14280 18776 14332 18785
rect 14556 18776 14608 18828
rect 15108 18776 15160 18828
rect 16764 18844 16816 18896
rect 17132 18844 17184 18896
rect 14004 18751 14056 18760
rect 14004 18717 14013 18751
rect 14013 18717 14047 18751
rect 14047 18717 14056 18751
rect 14004 18708 14056 18717
rect 16396 18819 16448 18828
rect 16396 18785 16405 18819
rect 16405 18785 16439 18819
rect 16439 18785 16448 18819
rect 16396 18776 16448 18785
rect 22284 18844 22336 18896
rect 11796 18640 11848 18649
rect 9772 18615 9824 18624
rect 9772 18581 9781 18615
rect 9781 18581 9815 18615
rect 9815 18581 9824 18615
rect 9772 18572 9824 18581
rect 13912 18615 13964 18624
rect 13912 18581 13921 18615
rect 13921 18581 13955 18615
rect 13955 18581 13964 18615
rect 13912 18572 13964 18581
rect 14188 18572 14240 18624
rect 19708 18776 19760 18828
rect 20352 18819 20404 18828
rect 20352 18785 20361 18819
rect 20361 18785 20395 18819
rect 20395 18785 20404 18819
rect 20352 18776 20404 18785
rect 20628 18776 20680 18828
rect 21088 18819 21140 18828
rect 21088 18785 21097 18819
rect 21097 18785 21131 18819
rect 21131 18785 21140 18819
rect 21088 18776 21140 18785
rect 22376 18776 22428 18828
rect 22928 18776 22980 18828
rect 21180 18708 21232 18760
rect 15292 18572 15344 18624
rect 15476 18615 15528 18624
rect 15476 18581 15485 18615
rect 15485 18581 15519 18615
rect 15519 18581 15528 18615
rect 15476 18572 15528 18581
rect 16488 18572 16540 18624
rect 17592 18572 17644 18624
rect 21364 18572 21416 18624
rect 22468 18572 22520 18624
rect 23020 18572 23072 18624
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 6552 18368 6604 18420
rect 14188 18368 14240 18420
rect 14280 18368 14332 18420
rect 16396 18368 16448 18420
rect 18420 18368 18472 18420
rect 5172 18300 5224 18352
rect 4160 18232 4212 18284
rect 4988 18232 5040 18284
rect 4620 18164 4672 18216
rect 4252 18139 4304 18148
rect 4252 18105 4261 18139
rect 4261 18105 4295 18139
rect 4295 18105 4304 18139
rect 4252 18096 4304 18105
rect 4344 18139 4396 18148
rect 4344 18105 4353 18139
rect 4353 18105 4387 18139
rect 4387 18105 4396 18139
rect 4896 18207 4948 18216
rect 4896 18173 4905 18207
rect 4905 18173 4939 18207
rect 4939 18173 4948 18207
rect 4896 18164 4948 18173
rect 5632 18207 5684 18216
rect 5632 18173 5641 18207
rect 5641 18173 5675 18207
rect 5675 18173 5684 18207
rect 5632 18164 5684 18173
rect 6092 18207 6144 18216
rect 6092 18173 6101 18207
rect 6101 18173 6135 18207
rect 6135 18173 6144 18207
rect 6092 18164 6144 18173
rect 8760 18300 8812 18352
rect 9036 18300 9088 18352
rect 10324 18232 10376 18284
rect 4344 18096 4396 18105
rect 5080 18096 5132 18148
rect 6000 18071 6052 18080
rect 6000 18037 6009 18071
rect 6009 18037 6043 18071
rect 6043 18037 6052 18071
rect 6000 18028 6052 18037
rect 6276 18028 6328 18080
rect 7012 18096 7064 18148
rect 7196 18096 7248 18148
rect 8484 18096 8536 18148
rect 9312 18164 9364 18216
rect 10048 18164 10100 18216
rect 10416 18164 10468 18216
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 11980 18275 12032 18284
rect 11980 18241 11989 18275
rect 11989 18241 12023 18275
rect 12023 18241 12032 18275
rect 11980 18232 12032 18241
rect 13912 18232 13964 18284
rect 14556 18232 14608 18284
rect 14648 18275 14700 18284
rect 14648 18241 14657 18275
rect 14657 18241 14691 18275
rect 14691 18241 14700 18275
rect 14648 18232 14700 18241
rect 15108 18232 15160 18284
rect 12072 18164 12124 18216
rect 14004 18164 14056 18216
rect 14740 18207 14792 18216
rect 14740 18173 14749 18207
rect 14749 18173 14783 18207
rect 14783 18173 14792 18207
rect 14740 18164 14792 18173
rect 14924 18207 14976 18216
rect 14924 18173 14933 18207
rect 14933 18173 14967 18207
rect 14967 18173 14976 18207
rect 14924 18164 14976 18173
rect 18144 18300 18196 18352
rect 21916 18368 21968 18420
rect 22008 18368 22060 18420
rect 22836 18368 22888 18420
rect 22928 18368 22980 18420
rect 17960 18275 18012 18284
rect 17960 18241 17969 18275
rect 17969 18241 18003 18275
rect 18003 18241 18012 18275
rect 17960 18232 18012 18241
rect 17592 18207 17644 18216
rect 17592 18173 17601 18207
rect 17601 18173 17635 18207
rect 17635 18173 17644 18207
rect 17592 18164 17644 18173
rect 17684 18207 17736 18216
rect 17684 18173 17693 18207
rect 17693 18173 17727 18207
rect 17727 18173 17736 18207
rect 17684 18164 17736 18173
rect 18236 18207 18288 18216
rect 18236 18173 18245 18207
rect 18245 18173 18279 18207
rect 18279 18173 18288 18207
rect 18236 18164 18288 18173
rect 18788 18207 18840 18216
rect 18788 18173 18797 18207
rect 18797 18173 18831 18207
rect 18831 18173 18840 18207
rect 18788 18164 18840 18173
rect 18972 18164 19024 18216
rect 19708 18207 19760 18216
rect 19708 18173 19717 18207
rect 19717 18173 19751 18207
rect 19751 18173 19760 18207
rect 19708 18164 19760 18173
rect 21364 18164 21416 18216
rect 21732 18164 21784 18216
rect 9496 18096 9548 18148
rect 12900 18096 12952 18148
rect 22744 18164 22796 18216
rect 21916 18139 21968 18148
rect 21916 18105 21950 18139
rect 21950 18105 21968 18139
rect 8760 18071 8812 18080
rect 8760 18037 8769 18071
rect 8769 18037 8803 18071
rect 8803 18037 8812 18071
rect 8760 18028 8812 18037
rect 8852 18071 8904 18080
rect 8852 18037 8861 18071
rect 8861 18037 8895 18071
rect 8895 18037 8904 18071
rect 8852 18028 8904 18037
rect 18604 18028 18656 18080
rect 21916 18096 21968 18105
rect 19892 18071 19944 18080
rect 19892 18037 19901 18071
rect 19901 18037 19935 18071
rect 19935 18037 19944 18071
rect 19892 18028 19944 18037
rect 22928 18028 22980 18080
rect 4322 17926 4374 17978
rect 4386 17926 4438 17978
rect 4450 17926 4502 17978
rect 4514 17926 4566 17978
rect 4578 17926 4630 17978
rect 4160 17824 4212 17876
rect 8760 17824 8812 17876
rect 9404 17824 9456 17876
rect 10048 17867 10100 17876
rect 10048 17833 10057 17867
rect 10057 17833 10091 17867
rect 10091 17833 10100 17867
rect 10048 17824 10100 17833
rect 18512 17824 18564 17876
rect 18604 17867 18656 17876
rect 18604 17833 18613 17867
rect 18613 17833 18647 17867
rect 18647 17833 18656 17867
rect 18604 17824 18656 17833
rect 22744 17867 22796 17876
rect 22744 17833 22753 17867
rect 22753 17833 22787 17867
rect 22787 17833 22796 17867
rect 22744 17824 22796 17833
rect 4804 17756 4856 17808
rect 4344 17731 4396 17740
rect 4344 17697 4353 17731
rect 4353 17697 4387 17731
rect 4387 17697 4396 17731
rect 4344 17688 4396 17697
rect 4620 17731 4672 17740
rect 4620 17697 4629 17731
rect 4629 17697 4663 17731
rect 4663 17697 4672 17731
rect 4620 17688 4672 17697
rect 5632 17756 5684 17808
rect 5908 17731 5960 17740
rect 4436 17663 4488 17672
rect 4436 17629 4445 17663
rect 4445 17629 4479 17663
rect 4479 17629 4488 17663
rect 4436 17620 4488 17629
rect 4896 17620 4948 17672
rect 5908 17697 5917 17731
rect 5917 17697 5951 17731
rect 5951 17697 5960 17731
rect 5908 17688 5960 17697
rect 7380 17731 7432 17740
rect 7380 17697 7389 17731
rect 7389 17697 7423 17731
rect 7423 17697 7432 17731
rect 7380 17688 7432 17697
rect 7472 17688 7524 17740
rect 9772 17756 9824 17808
rect 13912 17756 13964 17808
rect 9496 17688 9548 17740
rect 5632 17620 5684 17672
rect 6092 17552 6144 17604
rect 9220 17552 9272 17604
rect 14924 17688 14976 17740
rect 9864 17620 9916 17672
rect 16488 17731 16540 17740
rect 16488 17697 16497 17731
rect 16497 17697 16531 17731
rect 16531 17697 16540 17731
rect 16488 17688 16540 17697
rect 19892 17756 19944 17808
rect 16672 17688 16724 17740
rect 17224 17731 17276 17740
rect 17224 17697 17233 17731
rect 17233 17697 17267 17731
rect 17267 17697 17276 17731
rect 17224 17688 17276 17697
rect 16856 17620 16908 17672
rect 17592 17731 17644 17740
rect 17592 17697 17601 17731
rect 17601 17697 17635 17731
rect 17635 17697 17644 17731
rect 17592 17688 17644 17697
rect 17960 17688 18012 17740
rect 18144 17731 18196 17740
rect 18144 17697 18153 17731
rect 18153 17697 18187 17731
rect 18187 17697 18196 17731
rect 18144 17688 18196 17697
rect 18236 17688 18288 17740
rect 18696 17688 18748 17740
rect 19156 17688 19208 17740
rect 20904 17731 20956 17740
rect 20904 17697 20913 17731
rect 20913 17697 20947 17731
rect 20947 17697 20956 17731
rect 20904 17688 20956 17697
rect 22008 17688 22060 17740
rect 17132 17552 17184 17604
rect 21180 17620 21232 17672
rect 22836 17688 22888 17740
rect 23020 17731 23072 17740
rect 23020 17697 23029 17731
rect 23029 17697 23063 17731
rect 23063 17697 23072 17731
rect 23020 17688 23072 17697
rect 4712 17527 4764 17536
rect 4712 17493 4721 17527
rect 4721 17493 4755 17527
rect 4755 17493 4764 17527
rect 4712 17484 4764 17493
rect 8852 17484 8904 17536
rect 9864 17484 9916 17536
rect 16304 17484 16356 17536
rect 16764 17484 16816 17536
rect 18328 17527 18380 17536
rect 18328 17493 18337 17527
rect 18337 17493 18371 17527
rect 18371 17493 18380 17527
rect 18328 17484 18380 17493
rect 18788 17484 18840 17536
rect 20720 17527 20772 17536
rect 20720 17493 20729 17527
rect 20729 17493 20763 17527
rect 20763 17493 20772 17527
rect 20720 17484 20772 17493
rect 21548 17484 21600 17536
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 4252 17280 4304 17332
rect 4436 17076 4488 17128
rect 4712 17280 4764 17332
rect 5632 17323 5684 17332
rect 5632 17289 5641 17323
rect 5641 17289 5675 17323
rect 5675 17289 5684 17323
rect 5632 17280 5684 17289
rect 9496 17323 9548 17332
rect 9496 17289 9505 17323
rect 9505 17289 9539 17323
rect 9539 17289 9548 17323
rect 9496 17280 9548 17289
rect 13912 17323 13964 17332
rect 13912 17289 13921 17323
rect 13921 17289 13955 17323
rect 13955 17289 13964 17323
rect 13912 17280 13964 17289
rect 5540 17144 5592 17196
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 6276 17187 6328 17196
rect 6276 17153 6285 17187
rect 6285 17153 6319 17187
rect 6319 17153 6328 17187
rect 6276 17144 6328 17153
rect 7472 17212 7524 17264
rect 4988 17119 5040 17128
rect 4988 17085 4997 17119
rect 4997 17085 5031 17119
rect 5031 17085 5040 17119
rect 4988 17076 5040 17085
rect 6092 17076 6144 17128
rect 7380 17119 7432 17128
rect 7380 17085 7389 17119
rect 7389 17085 7423 17119
rect 7423 17085 7432 17119
rect 7380 17076 7432 17085
rect 8852 17119 8904 17128
rect 8852 17085 8861 17119
rect 8861 17085 8895 17119
rect 8895 17085 8904 17119
rect 8852 17076 8904 17085
rect 9220 17076 9272 17128
rect 9956 17076 10008 17128
rect 4344 17051 4396 17060
rect 4344 17017 4353 17051
rect 4353 17017 4387 17051
rect 4387 17017 4396 17051
rect 4344 17008 4396 17017
rect 5080 17008 5132 17060
rect 9036 17008 9088 17060
rect 10232 17119 10284 17128
rect 10232 17085 10241 17119
rect 10241 17085 10275 17119
rect 10275 17085 10284 17119
rect 10232 17076 10284 17085
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 11704 17119 11756 17128
rect 11704 17085 11713 17119
rect 11713 17085 11747 17119
rect 11747 17085 11756 17119
rect 11704 17076 11756 17085
rect 15660 17212 15712 17264
rect 16488 17280 16540 17332
rect 12900 17187 12952 17196
rect 12900 17153 12909 17187
rect 12909 17153 12943 17187
rect 12943 17153 12952 17187
rect 12900 17144 12952 17153
rect 14924 17187 14976 17196
rect 12900 17008 12952 17060
rect 4436 16940 4488 16992
rect 5172 16940 5224 16992
rect 8668 16983 8720 16992
rect 8668 16949 8677 16983
rect 8677 16949 8711 16983
rect 8711 16949 8720 16983
rect 8668 16940 8720 16949
rect 10232 16940 10284 16992
rect 10876 16940 10928 16992
rect 14924 17153 14933 17187
rect 14933 17153 14967 17187
rect 14967 17153 14976 17187
rect 14924 17144 14976 17153
rect 15476 17076 15528 17128
rect 15660 17076 15712 17128
rect 16304 17119 16356 17128
rect 16304 17085 16313 17119
rect 16313 17085 16347 17119
rect 16347 17085 16356 17119
rect 16304 17076 16356 17085
rect 16764 17119 16816 17128
rect 16764 17085 16773 17119
rect 16773 17085 16807 17119
rect 16807 17085 16816 17119
rect 16764 17076 16816 17085
rect 16856 17119 16908 17128
rect 16856 17085 16865 17119
rect 16865 17085 16899 17119
rect 16899 17085 16908 17119
rect 16856 17076 16908 17085
rect 17132 17323 17184 17332
rect 17132 17289 17141 17323
rect 17141 17289 17175 17323
rect 17175 17289 17184 17323
rect 17132 17280 17184 17289
rect 18236 17280 18288 17332
rect 18328 17323 18380 17332
rect 18328 17289 18337 17323
rect 18337 17289 18371 17323
rect 18371 17289 18380 17323
rect 18328 17280 18380 17289
rect 20904 17280 20956 17332
rect 21088 17280 21140 17332
rect 22008 17280 22060 17332
rect 17592 17144 17644 17196
rect 18420 17144 18472 17196
rect 17224 17119 17276 17128
rect 17224 17085 17233 17119
rect 17233 17085 17267 17119
rect 17267 17085 17276 17119
rect 17224 17076 17276 17085
rect 18052 17119 18104 17128
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 18052 17076 18104 17085
rect 18512 17119 18564 17128
rect 18512 17085 18521 17119
rect 18521 17085 18555 17119
rect 18555 17085 18564 17119
rect 18512 17076 18564 17085
rect 18696 17119 18748 17128
rect 18696 17085 18705 17119
rect 18705 17085 18739 17119
rect 18739 17085 18748 17119
rect 18696 17076 18748 17085
rect 15384 16983 15436 16992
rect 15384 16949 15393 16983
rect 15393 16949 15427 16983
rect 15427 16949 15436 16983
rect 15384 16940 15436 16949
rect 15568 16940 15620 16992
rect 16028 16940 16080 16992
rect 22744 17008 22796 17060
rect 19248 16940 19300 16992
rect 4322 16838 4374 16890
rect 4386 16838 4438 16890
rect 4450 16838 4502 16890
rect 4514 16838 4566 16890
rect 4578 16838 4630 16890
rect 4252 16779 4304 16788
rect 4252 16745 4261 16779
rect 4261 16745 4295 16779
rect 4295 16745 4304 16779
rect 4252 16736 4304 16745
rect 4068 16668 4120 16720
rect 4712 16668 4764 16720
rect 5448 16736 5500 16788
rect 9036 16779 9088 16788
rect 9036 16745 9045 16779
rect 9045 16745 9079 16779
rect 9079 16745 9088 16779
rect 9036 16736 9088 16745
rect 9496 16736 9548 16788
rect 4160 16643 4212 16652
rect 4160 16609 4169 16643
rect 4169 16609 4203 16643
rect 4203 16609 4212 16643
rect 4160 16600 4212 16609
rect 5172 16643 5224 16652
rect 5172 16609 5181 16643
rect 5181 16609 5215 16643
rect 5215 16609 5224 16643
rect 5172 16600 5224 16609
rect 4252 16532 4304 16584
rect 4712 16575 4764 16584
rect 4712 16541 4721 16575
rect 4721 16541 4755 16575
rect 4755 16541 4764 16575
rect 4712 16532 4764 16541
rect 6276 16600 6328 16652
rect 7564 16600 7616 16652
rect 8852 16643 8904 16652
rect 8852 16609 8861 16643
rect 8861 16609 8895 16643
rect 8895 16609 8904 16643
rect 8852 16600 8904 16609
rect 9404 16711 9456 16720
rect 9404 16677 9413 16711
rect 9413 16677 9447 16711
rect 9447 16677 9456 16711
rect 9404 16668 9456 16677
rect 9220 16600 9272 16652
rect 13544 16736 13596 16788
rect 14556 16779 14608 16788
rect 14556 16745 14565 16779
rect 14565 16745 14599 16779
rect 14599 16745 14608 16779
rect 14556 16736 14608 16745
rect 15660 16736 15712 16788
rect 13360 16643 13412 16652
rect 13360 16609 13369 16643
rect 13369 16609 13403 16643
rect 13403 16609 13412 16643
rect 13360 16600 13412 16609
rect 13544 16643 13596 16652
rect 13544 16609 13553 16643
rect 13553 16609 13587 16643
rect 13587 16609 13596 16643
rect 13544 16600 13596 16609
rect 14188 16668 14240 16720
rect 13728 16643 13780 16652
rect 13728 16609 13737 16643
rect 13737 16609 13771 16643
rect 13771 16609 13780 16643
rect 13728 16600 13780 16609
rect 14280 16643 14332 16652
rect 14280 16609 14289 16643
rect 14289 16609 14323 16643
rect 14323 16609 14332 16643
rect 14280 16600 14332 16609
rect 16028 16668 16080 16720
rect 17132 16736 17184 16788
rect 18512 16736 18564 16788
rect 16672 16711 16724 16720
rect 16672 16677 16681 16711
rect 16681 16677 16715 16711
rect 16715 16677 16724 16711
rect 16672 16668 16724 16677
rect 14464 16600 14516 16652
rect 15016 16643 15068 16652
rect 15016 16609 15025 16643
rect 15025 16609 15059 16643
rect 15059 16609 15068 16643
rect 15016 16600 15068 16609
rect 15200 16643 15252 16652
rect 15200 16609 15209 16643
rect 15209 16609 15243 16643
rect 15243 16609 15252 16643
rect 15200 16600 15252 16609
rect 15384 16600 15436 16652
rect 15108 16532 15160 16584
rect 15660 16532 15712 16584
rect 16396 16532 16448 16584
rect 18696 16600 18748 16652
rect 19708 16668 19760 16720
rect 21824 16711 21876 16720
rect 21824 16677 21833 16711
rect 21833 16677 21867 16711
rect 21867 16677 21876 16711
rect 21824 16668 21876 16677
rect 19248 16600 19300 16652
rect 21548 16643 21600 16652
rect 21548 16609 21557 16643
rect 21557 16609 21591 16643
rect 21591 16609 21600 16643
rect 21548 16600 21600 16609
rect 22100 16532 22152 16584
rect 22560 16532 22612 16584
rect 5080 16464 5132 16516
rect 10232 16464 10284 16516
rect 15568 16464 15620 16516
rect 16212 16464 16264 16516
rect 18052 16464 18104 16516
rect 5356 16439 5408 16448
rect 5356 16405 5365 16439
rect 5365 16405 5399 16439
rect 5399 16405 5408 16439
rect 5356 16396 5408 16405
rect 9680 16396 9732 16448
rect 9772 16439 9824 16448
rect 9772 16405 9781 16439
rect 9781 16405 9815 16439
rect 9815 16405 9824 16439
rect 9772 16396 9824 16405
rect 15384 16439 15436 16448
rect 15384 16405 15393 16439
rect 15393 16405 15427 16439
rect 15427 16405 15436 16439
rect 15384 16396 15436 16405
rect 16304 16439 16356 16448
rect 16304 16405 16313 16439
rect 16313 16405 16347 16439
rect 16347 16405 16356 16439
rect 16304 16396 16356 16405
rect 21640 16439 21692 16448
rect 21640 16405 21649 16439
rect 21649 16405 21683 16439
rect 21683 16405 21692 16439
rect 21640 16396 21692 16405
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 13728 16192 13780 16244
rect 15108 16192 15160 16244
rect 16304 16192 16356 16244
rect 7104 16124 7156 16176
rect 5356 16099 5408 16108
rect 5356 16065 5365 16099
rect 5365 16065 5399 16099
rect 5399 16065 5408 16099
rect 5356 16056 5408 16065
rect 6736 16056 6788 16108
rect 5264 16031 5316 16040
rect 5264 15997 5273 16031
rect 5273 15997 5307 16031
rect 5307 15997 5316 16031
rect 5264 15988 5316 15997
rect 7012 15988 7064 16040
rect 6920 15963 6972 15972
rect 6920 15929 6929 15963
rect 6929 15929 6963 15963
rect 6963 15929 6972 15963
rect 6920 15920 6972 15929
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 8024 15920 8076 15972
rect 11612 16056 11664 16108
rect 11428 15988 11480 16040
rect 13544 16124 13596 16176
rect 13360 16056 13412 16108
rect 15200 16124 15252 16176
rect 16764 16192 16816 16244
rect 18604 16192 18656 16244
rect 19432 16192 19484 16244
rect 21548 16192 21600 16244
rect 22100 16192 22152 16244
rect 22652 16192 22704 16244
rect 13452 15988 13504 16040
rect 15108 16056 15160 16108
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 15016 15988 15068 16040
rect 15200 16031 15252 16040
rect 15200 15997 15209 16031
rect 15209 15997 15243 16031
rect 15243 15997 15252 16031
rect 15200 15988 15252 15997
rect 15660 16056 15712 16108
rect 16672 16124 16724 16176
rect 16948 16167 17000 16176
rect 16948 16133 16957 16167
rect 16957 16133 16991 16167
rect 16991 16133 17000 16167
rect 16948 16124 17000 16133
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 16304 16099 16356 16108
rect 16304 16065 16313 16099
rect 16313 16065 16347 16099
rect 16347 16065 16356 16099
rect 16304 16056 16356 16065
rect 19524 16124 19576 16176
rect 19708 16124 19760 16176
rect 16488 15988 16540 16040
rect 16764 16031 16816 16040
rect 16764 15997 16773 16031
rect 16773 15997 16807 16031
rect 16807 15997 16816 16031
rect 16764 15988 16816 15997
rect 19432 16056 19484 16108
rect 19156 16031 19208 16040
rect 19156 15997 19165 16031
rect 19165 15997 19199 16031
rect 19199 15997 19208 16031
rect 19156 15988 19208 15997
rect 19248 16031 19300 16040
rect 19248 15997 19257 16031
rect 19257 15997 19291 16031
rect 19291 15997 19300 16031
rect 19248 15988 19300 15997
rect 20352 15988 20404 16040
rect 21456 16056 21508 16108
rect 22192 16056 22244 16108
rect 21640 16031 21692 16040
rect 12992 15963 13044 15972
rect 12992 15929 13001 15963
rect 13001 15929 13035 15963
rect 13035 15929 13044 15963
rect 12992 15920 13044 15929
rect 11428 15852 11480 15904
rect 11704 15852 11756 15904
rect 13544 15852 13596 15904
rect 14280 15895 14332 15904
rect 14280 15861 14289 15895
rect 14289 15861 14323 15895
rect 14323 15861 14332 15895
rect 14280 15852 14332 15861
rect 15384 15852 15436 15904
rect 16304 15852 16356 15904
rect 16580 15895 16632 15904
rect 16580 15861 16589 15895
rect 16589 15861 16623 15895
rect 16623 15861 16632 15895
rect 16580 15852 16632 15861
rect 16672 15852 16724 15904
rect 19524 15895 19576 15904
rect 19524 15861 19533 15895
rect 19533 15861 19567 15895
rect 19567 15861 19576 15895
rect 19524 15852 19576 15861
rect 19708 15852 19760 15904
rect 20812 15920 20864 15972
rect 21640 15997 21649 16031
rect 21649 15997 21683 16031
rect 21683 15997 21692 16031
rect 21640 15988 21692 15997
rect 20720 15895 20772 15904
rect 20720 15861 20729 15895
rect 20729 15861 20763 15895
rect 20763 15861 20772 15895
rect 20720 15852 20772 15861
rect 21640 15852 21692 15904
rect 4322 15750 4374 15802
rect 4386 15750 4438 15802
rect 4450 15750 4502 15802
rect 4514 15750 4566 15802
rect 4578 15750 4630 15802
rect 4252 15648 4304 15700
rect 4804 15648 4856 15700
rect 15200 15648 15252 15700
rect 20168 15648 20220 15700
rect 20812 15691 20864 15700
rect 20812 15657 20821 15691
rect 20821 15657 20855 15691
rect 20855 15657 20864 15691
rect 20812 15648 20864 15657
rect 4068 15555 4120 15564
rect 4068 15521 4077 15555
rect 4077 15521 4111 15555
rect 4111 15521 4120 15555
rect 4068 15512 4120 15521
rect 5080 15512 5132 15564
rect 5816 15512 5868 15564
rect 6000 15555 6052 15564
rect 6000 15521 6009 15555
rect 6009 15521 6043 15555
rect 6043 15521 6052 15555
rect 6000 15512 6052 15521
rect 7564 15512 7616 15564
rect 4712 15444 4764 15496
rect 6092 15487 6144 15496
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 7196 15487 7248 15496
rect 6000 15376 6052 15428
rect 7196 15453 7205 15487
rect 7205 15453 7239 15487
rect 7239 15453 7248 15487
rect 7196 15444 7248 15453
rect 8668 15444 8720 15496
rect 10140 15580 10192 15632
rect 11520 15580 11572 15632
rect 16488 15623 16540 15632
rect 16488 15589 16497 15623
rect 16497 15589 16531 15623
rect 16531 15589 16540 15623
rect 16488 15580 16540 15589
rect 16580 15580 16632 15632
rect 11428 15512 11480 15564
rect 12992 15555 13044 15564
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 13452 15512 13504 15564
rect 16212 15512 16264 15564
rect 7012 15419 7064 15428
rect 7012 15385 7021 15419
rect 7021 15385 7055 15419
rect 7055 15385 7064 15419
rect 7012 15376 7064 15385
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 13820 15444 13872 15496
rect 16672 15555 16724 15564
rect 16672 15521 16681 15555
rect 16681 15521 16715 15555
rect 16715 15521 16724 15555
rect 16672 15512 16724 15521
rect 16948 15555 17000 15564
rect 16948 15521 16957 15555
rect 16957 15521 16991 15555
rect 16991 15521 17000 15555
rect 16948 15512 17000 15521
rect 17316 15555 17368 15564
rect 17316 15521 17325 15555
rect 17325 15521 17359 15555
rect 17359 15521 17368 15555
rect 17316 15512 17368 15521
rect 19524 15555 19576 15564
rect 19524 15521 19533 15555
rect 19533 15521 19567 15555
rect 19567 15521 19576 15555
rect 19524 15512 19576 15521
rect 19708 15555 19760 15564
rect 19708 15521 19717 15555
rect 19717 15521 19751 15555
rect 19751 15521 19760 15555
rect 19708 15512 19760 15521
rect 16856 15444 16908 15496
rect 20720 15555 20772 15564
rect 20720 15521 20729 15555
rect 20729 15521 20763 15555
rect 20763 15521 20772 15555
rect 20720 15512 20772 15521
rect 22192 15512 22244 15564
rect 9680 15376 9732 15428
rect 12072 15419 12124 15428
rect 12072 15385 12081 15419
rect 12081 15385 12115 15419
rect 12115 15385 12124 15419
rect 12072 15376 12124 15385
rect 9956 15308 10008 15360
rect 10048 15308 10100 15360
rect 15936 15308 15988 15360
rect 16764 15351 16816 15360
rect 16764 15317 16773 15351
rect 16773 15317 16807 15351
rect 16807 15317 16816 15351
rect 16764 15308 16816 15317
rect 17132 15308 17184 15360
rect 18788 15308 18840 15360
rect 19708 15308 19760 15360
rect 20812 15376 20864 15428
rect 20536 15308 20588 15360
rect 20720 15308 20772 15360
rect 21640 15487 21692 15496
rect 21640 15453 21649 15487
rect 21649 15453 21683 15487
rect 21683 15453 21692 15487
rect 21640 15444 21692 15453
rect 20996 15351 21048 15360
rect 20996 15317 21005 15351
rect 21005 15317 21039 15351
rect 21039 15317 21048 15351
rect 20996 15308 21048 15317
rect 22100 15351 22152 15360
rect 22100 15317 22109 15351
rect 22109 15317 22143 15351
rect 22143 15317 22152 15351
rect 22100 15308 22152 15317
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 4160 15104 4212 15156
rect 4804 14943 4856 14952
rect 4804 14909 4813 14943
rect 4813 14909 4847 14943
rect 4847 14909 4856 14943
rect 4804 14900 4856 14909
rect 5172 14900 5224 14952
rect 6920 15104 6972 15156
rect 7196 15104 7248 15156
rect 11888 15104 11940 15156
rect 6000 15036 6052 15088
rect 6092 15011 6144 15020
rect 6092 14977 6101 15011
rect 6101 14977 6135 15011
rect 6135 14977 6144 15011
rect 6092 14968 6144 14977
rect 5448 14900 5500 14952
rect 7104 14968 7156 15020
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 7012 14943 7064 14952
rect 7012 14909 7022 14943
rect 7022 14909 7056 14943
rect 7056 14909 7064 14943
rect 7012 14900 7064 14909
rect 10140 14900 10192 14952
rect 11244 14900 11296 14952
rect 14280 15104 14332 15156
rect 12808 15036 12860 15088
rect 16856 15104 16908 15156
rect 17040 15147 17092 15156
rect 17040 15113 17049 15147
rect 17049 15113 17083 15147
rect 17083 15113 17092 15147
rect 17040 15104 17092 15113
rect 18696 15104 18748 15156
rect 20996 15104 21048 15156
rect 11520 14943 11572 14952
rect 11520 14909 11529 14943
rect 11529 14909 11563 14943
rect 11563 14909 11572 14943
rect 11520 14900 11572 14909
rect 18604 14968 18656 15020
rect 19156 15011 19208 15020
rect 12072 14900 12124 14952
rect 4252 14764 4304 14816
rect 5632 14764 5684 14816
rect 6920 14764 6972 14816
rect 9680 14764 9732 14816
rect 10324 14764 10376 14816
rect 13544 14943 13596 14952
rect 13544 14909 13553 14943
rect 13553 14909 13587 14943
rect 13587 14909 13596 14943
rect 13544 14900 13596 14909
rect 13728 14900 13780 14952
rect 15936 14943 15988 14952
rect 15936 14909 15970 14943
rect 15970 14909 15988 14943
rect 12164 14764 12216 14816
rect 13176 14764 13228 14816
rect 13728 14764 13780 14816
rect 15936 14900 15988 14909
rect 17316 14900 17368 14952
rect 17960 14943 18012 14952
rect 17960 14909 17969 14943
rect 17969 14909 18003 14943
rect 18003 14909 18012 14943
rect 17960 14900 18012 14909
rect 18052 14943 18104 14952
rect 18052 14909 18061 14943
rect 18061 14909 18095 14943
rect 18095 14909 18104 14943
rect 19156 14977 19165 15011
rect 19165 14977 19199 15011
rect 19199 14977 19208 15011
rect 19156 14968 19208 14977
rect 19708 15011 19760 15020
rect 19708 14977 19717 15011
rect 19717 14977 19751 15011
rect 19751 14977 19760 15011
rect 19708 14968 19760 14977
rect 20904 14968 20956 15020
rect 21456 15011 21508 15020
rect 21456 14977 21465 15011
rect 21465 14977 21499 15011
rect 21499 14977 21508 15011
rect 21456 14968 21508 14977
rect 18052 14900 18104 14909
rect 19248 14900 19300 14952
rect 20444 14900 20496 14952
rect 20536 14943 20588 14952
rect 20536 14909 20545 14943
rect 20545 14909 20579 14943
rect 20579 14909 20588 14943
rect 20536 14900 20588 14909
rect 21364 14943 21416 14952
rect 21364 14909 21373 14943
rect 21373 14909 21407 14943
rect 21407 14909 21416 14943
rect 21364 14900 21416 14909
rect 22100 14900 22152 14952
rect 22652 14943 22704 14952
rect 22652 14909 22661 14943
rect 22661 14909 22695 14943
rect 22695 14909 22704 14943
rect 22652 14900 22704 14909
rect 16396 14832 16448 14884
rect 17776 14832 17828 14884
rect 18328 14832 18380 14884
rect 19432 14832 19484 14884
rect 15936 14764 15988 14816
rect 22376 14807 22428 14816
rect 22376 14773 22385 14807
rect 22385 14773 22419 14807
rect 22419 14773 22428 14807
rect 22376 14764 22428 14773
rect 4322 14662 4374 14714
rect 4386 14662 4438 14714
rect 4450 14662 4502 14714
rect 4514 14662 4566 14714
rect 4578 14662 4630 14714
rect 9956 14560 10008 14612
rect 4252 14492 4304 14544
rect 8024 14492 8076 14544
rect 7196 14424 7248 14476
rect 8300 14467 8352 14476
rect 8300 14433 8309 14467
rect 8309 14433 8343 14467
rect 8343 14433 8352 14467
rect 8300 14424 8352 14433
rect 8116 14356 8168 14408
rect 9220 14424 9272 14476
rect 9680 14492 9732 14544
rect 10232 14492 10284 14544
rect 10324 14535 10376 14544
rect 10324 14501 10333 14535
rect 10333 14501 10367 14535
rect 10367 14501 10376 14535
rect 10600 14535 10652 14544
rect 10324 14492 10376 14501
rect 10600 14501 10611 14535
rect 10611 14501 10652 14535
rect 10600 14492 10652 14501
rect 11428 14560 11480 14612
rect 14464 14560 14516 14612
rect 17316 14560 17368 14612
rect 9588 14356 9640 14408
rect 9864 14424 9916 14476
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 8944 14288 8996 14340
rect 9864 14288 9916 14340
rect 5632 14263 5684 14272
rect 5632 14229 5641 14263
rect 5641 14229 5675 14263
rect 5675 14229 5684 14263
rect 5632 14220 5684 14229
rect 8392 14220 8444 14272
rect 9772 14220 9824 14272
rect 9956 14263 10008 14272
rect 9956 14229 9965 14263
rect 9965 14229 9999 14263
rect 9999 14229 10008 14263
rect 9956 14220 10008 14229
rect 10140 14220 10192 14272
rect 10416 14263 10468 14272
rect 10416 14229 10425 14263
rect 10425 14229 10459 14263
rect 10459 14229 10468 14263
rect 10416 14220 10468 14229
rect 10692 14356 10744 14408
rect 12072 14424 12124 14476
rect 16764 14492 16816 14544
rect 13176 14467 13228 14476
rect 13176 14433 13185 14467
rect 13185 14433 13219 14467
rect 13219 14433 13228 14467
rect 13176 14424 13228 14433
rect 13544 14424 13596 14476
rect 13728 14467 13780 14476
rect 13728 14433 13737 14467
rect 13737 14433 13771 14467
rect 13771 14433 13780 14467
rect 13728 14424 13780 14433
rect 13912 14424 13964 14476
rect 17960 14560 18012 14612
rect 19432 14603 19484 14612
rect 19432 14569 19441 14603
rect 19441 14569 19475 14603
rect 19475 14569 19484 14603
rect 19432 14560 19484 14569
rect 18328 14492 18380 14544
rect 17776 14467 17828 14476
rect 17776 14433 17785 14467
rect 17785 14433 17819 14467
rect 17819 14433 17828 14467
rect 17776 14424 17828 14433
rect 18512 14467 18564 14476
rect 18512 14433 18521 14467
rect 18521 14433 18555 14467
rect 18555 14433 18564 14467
rect 18512 14424 18564 14433
rect 18972 14467 19024 14476
rect 18972 14433 18981 14467
rect 18981 14433 19015 14467
rect 19015 14433 19024 14467
rect 18972 14424 19024 14433
rect 21824 14560 21876 14612
rect 22836 14560 22888 14612
rect 13268 14399 13320 14408
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 13268 14356 13320 14365
rect 15936 14356 15988 14408
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 18788 14356 18840 14408
rect 21732 14424 21784 14476
rect 21824 14467 21876 14476
rect 21824 14433 21833 14467
rect 21833 14433 21867 14467
rect 21867 14433 21876 14467
rect 21824 14424 21876 14433
rect 21640 14356 21692 14408
rect 22008 14467 22060 14476
rect 22008 14433 22017 14467
rect 22017 14433 22051 14467
rect 22051 14433 22060 14467
rect 22008 14424 22060 14433
rect 22192 14424 22244 14476
rect 22468 14424 22520 14476
rect 22284 14399 22336 14408
rect 22284 14365 22293 14399
rect 22293 14365 22327 14399
rect 22327 14365 22336 14399
rect 22284 14356 22336 14365
rect 22560 14356 22612 14408
rect 12716 14220 12768 14272
rect 13820 14220 13872 14272
rect 18052 14263 18104 14272
rect 18052 14229 18061 14263
rect 18061 14229 18095 14263
rect 18095 14229 18104 14263
rect 18052 14220 18104 14229
rect 18236 14263 18288 14272
rect 18236 14229 18245 14263
rect 18245 14229 18279 14263
rect 18279 14229 18288 14263
rect 18236 14220 18288 14229
rect 19064 14263 19116 14272
rect 19064 14229 19073 14263
rect 19073 14229 19107 14263
rect 19107 14229 19116 14263
rect 19064 14220 19116 14229
rect 22376 14220 22428 14272
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 5172 14016 5224 14068
rect 9036 14016 9088 14068
rect 9588 14059 9640 14068
rect 9588 14025 9597 14059
rect 9597 14025 9631 14059
rect 9631 14025 9640 14059
rect 9588 14016 9640 14025
rect 9220 13948 9272 14000
rect 10416 14016 10468 14068
rect 12440 14016 12492 14068
rect 6920 13880 6972 13932
rect 8116 13880 8168 13932
rect 8944 13880 8996 13932
rect 7196 13812 7248 13864
rect 8392 13855 8444 13864
rect 8392 13821 8401 13855
rect 8401 13821 8435 13855
rect 8435 13821 8444 13855
rect 8392 13812 8444 13821
rect 8576 13855 8628 13864
rect 8576 13821 8585 13855
rect 8585 13821 8619 13855
rect 8619 13821 8628 13855
rect 8576 13812 8628 13821
rect 8760 13812 8812 13864
rect 5448 13744 5500 13796
rect 9036 13812 9088 13864
rect 9772 13880 9824 13932
rect 12532 13948 12584 14000
rect 9864 13812 9916 13864
rect 10140 13812 10192 13864
rect 10324 13855 10376 13864
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 12440 13880 12492 13932
rect 13820 14059 13872 14068
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 16764 14016 16816 14068
rect 12716 13923 12768 13932
rect 12716 13889 12725 13923
rect 12725 13889 12759 13923
rect 12759 13889 12768 13923
rect 12716 13880 12768 13889
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 8760 13719 8812 13728
rect 8760 13685 8769 13719
rect 8769 13685 8803 13719
rect 8803 13685 8812 13719
rect 8760 13676 8812 13685
rect 9588 13744 9640 13796
rect 10140 13676 10192 13728
rect 11060 13812 11112 13864
rect 11428 13855 11480 13864
rect 11428 13821 11437 13855
rect 11437 13821 11471 13855
rect 11471 13821 11480 13855
rect 11428 13812 11480 13821
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 13820 13880 13872 13932
rect 10416 13676 10468 13728
rect 11060 13676 11112 13728
rect 11152 13719 11204 13728
rect 11152 13685 11161 13719
rect 11161 13685 11195 13719
rect 11195 13685 11204 13719
rect 11152 13676 11204 13685
rect 13176 13812 13228 13864
rect 13544 13812 13596 13864
rect 14096 13948 14148 14000
rect 18052 14016 18104 14068
rect 19064 14059 19116 14068
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 17776 13948 17828 14000
rect 17960 13991 18012 14000
rect 17960 13957 17969 13991
rect 17969 13957 18003 13991
rect 18003 13957 18012 13991
rect 17960 13948 18012 13957
rect 14372 13923 14424 13932
rect 14372 13889 14381 13923
rect 14381 13889 14415 13923
rect 14415 13889 14424 13923
rect 14372 13880 14424 13889
rect 17132 13880 17184 13932
rect 21272 14016 21324 14068
rect 21548 14016 21600 14068
rect 12624 13744 12676 13796
rect 13636 13787 13688 13796
rect 13636 13753 13645 13787
rect 13645 13753 13679 13787
rect 13679 13753 13688 13787
rect 13636 13744 13688 13753
rect 15292 13812 15344 13864
rect 15476 13744 15528 13796
rect 17224 13787 17276 13796
rect 17224 13753 17233 13787
rect 17233 13753 17267 13787
rect 17267 13753 17276 13787
rect 17224 13744 17276 13753
rect 12808 13676 12860 13728
rect 16028 13719 16080 13728
rect 16028 13685 16037 13719
rect 16037 13685 16071 13719
rect 16071 13685 16080 13719
rect 16028 13676 16080 13685
rect 17132 13676 17184 13728
rect 17776 13855 17828 13864
rect 17776 13821 17785 13855
rect 17785 13821 17819 13855
rect 17819 13821 17828 13855
rect 17776 13812 17828 13821
rect 22836 13948 22888 14000
rect 18236 13812 18288 13864
rect 20904 13812 20956 13864
rect 22744 13880 22796 13932
rect 18696 13787 18748 13796
rect 18696 13753 18705 13787
rect 18705 13753 18739 13787
rect 18739 13753 18748 13787
rect 18696 13744 18748 13753
rect 21364 13676 21416 13728
rect 21824 13719 21876 13728
rect 21824 13685 21833 13719
rect 21833 13685 21867 13719
rect 21867 13685 21876 13719
rect 21824 13676 21876 13685
rect 4322 13574 4374 13626
rect 4386 13574 4438 13626
rect 4450 13574 4502 13626
rect 4514 13574 4566 13626
rect 4578 13574 4630 13626
rect 5356 13515 5408 13524
rect 5356 13481 5365 13515
rect 5365 13481 5399 13515
rect 5399 13481 5408 13515
rect 5356 13472 5408 13481
rect 6368 13472 6420 13524
rect 8392 13472 8444 13524
rect 10416 13515 10468 13524
rect 10416 13481 10425 13515
rect 10425 13481 10459 13515
rect 10459 13481 10468 13515
rect 10416 13472 10468 13481
rect 12716 13472 12768 13524
rect 12808 13515 12860 13524
rect 12808 13481 12817 13515
rect 12817 13481 12851 13515
rect 12851 13481 12860 13515
rect 12808 13472 12860 13481
rect 13728 13472 13780 13524
rect 15476 13472 15528 13524
rect 16764 13515 16816 13524
rect 16764 13481 16773 13515
rect 16773 13481 16807 13515
rect 16807 13481 16816 13515
rect 16764 13472 16816 13481
rect 17132 13515 17184 13524
rect 17132 13481 17141 13515
rect 17141 13481 17175 13515
rect 17175 13481 17184 13515
rect 17132 13472 17184 13481
rect 18788 13472 18840 13524
rect 21732 13472 21784 13524
rect 8116 13447 8168 13456
rect 8116 13413 8125 13447
rect 8125 13413 8159 13447
rect 8159 13413 8168 13447
rect 8116 13404 8168 13413
rect 8484 13404 8536 13456
rect 8760 13447 8812 13456
rect 8760 13413 8769 13447
rect 8769 13413 8803 13447
rect 8803 13413 8812 13447
rect 8760 13404 8812 13413
rect 5264 13379 5316 13388
rect 5264 13345 5273 13379
rect 5273 13345 5307 13379
rect 5307 13345 5316 13379
rect 5264 13336 5316 13345
rect 6184 13379 6236 13388
rect 6184 13345 6193 13379
rect 6193 13345 6227 13379
rect 6227 13345 6236 13379
rect 6184 13336 6236 13345
rect 8576 13336 8628 13388
rect 8944 13379 8996 13388
rect 8944 13345 8953 13379
rect 8953 13345 8987 13379
rect 8987 13345 8996 13379
rect 8944 13336 8996 13345
rect 6828 13268 6880 13320
rect 9956 13379 10008 13388
rect 9956 13345 9965 13379
rect 9965 13345 9999 13379
rect 9999 13345 10008 13379
rect 9956 13336 10008 13345
rect 12532 13404 12584 13456
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 10048 13268 10100 13320
rect 12348 13379 12400 13388
rect 12348 13345 12357 13379
rect 12357 13345 12391 13379
rect 12391 13345 12400 13379
rect 12348 13336 12400 13345
rect 12624 13379 12676 13388
rect 12624 13345 12633 13379
rect 12633 13345 12667 13379
rect 12667 13345 12676 13379
rect 12624 13336 12676 13345
rect 13268 13379 13320 13388
rect 13268 13345 13281 13379
rect 13281 13345 13320 13379
rect 13268 13336 13320 13345
rect 13820 13379 13872 13388
rect 13820 13345 13829 13379
rect 13829 13345 13863 13379
rect 13863 13345 13872 13379
rect 13820 13336 13872 13345
rect 14372 13336 14424 13388
rect 16028 13404 16080 13456
rect 14004 13311 14056 13320
rect 14004 13277 14013 13311
rect 14013 13277 14047 13311
rect 14047 13277 14056 13311
rect 14004 13268 14056 13277
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16396 13379 16448 13388
rect 16396 13345 16405 13379
rect 16405 13345 16439 13379
rect 16439 13345 16448 13379
rect 18052 13404 18104 13456
rect 16396 13336 16448 13345
rect 16304 13268 16356 13320
rect 17868 13336 17920 13388
rect 18420 13447 18472 13456
rect 18420 13413 18445 13447
rect 18445 13413 18472 13447
rect 18420 13404 18472 13413
rect 18328 13336 18380 13388
rect 19156 13336 19208 13388
rect 17040 13268 17092 13320
rect 18052 13268 18104 13320
rect 20812 13404 20864 13456
rect 22100 13404 22152 13456
rect 21364 13336 21416 13388
rect 21640 13336 21692 13388
rect 22008 13379 22060 13388
rect 22008 13345 22017 13379
rect 22017 13345 22051 13379
rect 22051 13345 22060 13379
rect 22008 13336 22060 13345
rect 22652 13379 22704 13388
rect 22652 13345 22661 13379
rect 22661 13345 22695 13379
rect 22695 13345 22704 13379
rect 22652 13336 22704 13345
rect 20444 13311 20496 13320
rect 20444 13277 20453 13311
rect 20453 13277 20487 13311
rect 20487 13277 20496 13311
rect 20444 13268 20496 13277
rect 20536 13311 20588 13320
rect 20536 13277 20545 13311
rect 20545 13277 20579 13311
rect 20579 13277 20588 13311
rect 20536 13268 20588 13277
rect 20628 13311 20680 13320
rect 20628 13277 20637 13311
rect 20637 13277 20671 13311
rect 20671 13277 20680 13311
rect 20628 13268 20680 13277
rect 4896 13175 4948 13184
rect 4896 13141 4905 13175
rect 4905 13141 4939 13175
rect 4939 13141 4948 13175
rect 4896 13132 4948 13141
rect 5816 13175 5868 13184
rect 5816 13141 5825 13175
rect 5825 13141 5859 13175
rect 5859 13141 5868 13175
rect 5816 13132 5868 13141
rect 8208 13132 8260 13184
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 9772 13175 9824 13184
rect 9772 13141 9781 13175
rect 9781 13141 9815 13175
rect 9815 13141 9824 13175
rect 9772 13132 9824 13141
rect 13636 13132 13688 13184
rect 19340 13200 19392 13252
rect 18512 13132 18564 13184
rect 19708 13132 19760 13184
rect 19800 13175 19852 13184
rect 19800 13141 19809 13175
rect 19809 13141 19843 13175
rect 19843 13141 19852 13175
rect 19800 13132 19852 13141
rect 20996 13200 21048 13252
rect 21272 13200 21324 13252
rect 20628 13132 20680 13184
rect 21088 13132 21140 13184
rect 21916 13175 21968 13184
rect 21916 13141 21925 13175
rect 21925 13141 21959 13175
rect 21959 13141 21968 13175
rect 21916 13132 21968 13141
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 5908 12971 5960 12980
rect 5908 12937 5917 12971
rect 5917 12937 5951 12971
rect 5951 12937 5960 12971
rect 5908 12928 5960 12937
rect 6184 12928 6236 12980
rect 11060 12928 11112 12980
rect 9036 12792 9088 12844
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 12348 12928 12400 12980
rect 12440 12971 12492 12980
rect 12440 12937 12449 12971
rect 12449 12937 12483 12971
rect 12483 12937 12492 12971
rect 12440 12928 12492 12937
rect 15200 12928 15252 12980
rect 20444 12928 20496 12980
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 21088 12971 21140 12980
rect 21088 12937 21097 12971
rect 21097 12937 21131 12971
rect 21131 12937 21140 12971
rect 21088 12928 21140 12937
rect 21364 12928 21416 12980
rect 4252 12656 4304 12708
rect 5816 12724 5868 12776
rect 5448 12656 5500 12708
rect 8392 12724 8444 12776
rect 9128 12767 9180 12776
rect 9128 12733 9137 12767
rect 9137 12733 9171 12767
rect 9171 12733 9180 12767
rect 9128 12724 9180 12733
rect 9312 12767 9364 12776
rect 9312 12733 9321 12767
rect 9321 12733 9355 12767
rect 9355 12733 9364 12767
rect 9312 12724 9364 12733
rect 18420 12860 18472 12912
rect 6460 12656 6512 12708
rect 6828 12656 6880 12708
rect 7380 12631 7432 12640
rect 7380 12597 7389 12631
rect 7389 12597 7423 12631
rect 7423 12597 7432 12631
rect 7380 12588 7432 12597
rect 9680 12656 9732 12708
rect 11428 12767 11480 12776
rect 11428 12733 11437 12767
rect 11437 12733 11471 12767
rect 11471 12733 11480 12767
rect 11428 12724 11480 12733
rect 11980 12767 12032 12776
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 12532 12767 12584 12776
rect 12532 12733 12541 12767
rect 12541 12733 12575 12767
rect 12575 12733 12584 12767
rect 12532 12724 12584 12733
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 13636 12724 13688 12776
rect 11520 12656 11572 12708
rect 12900 12656 12952 12708
rect 18052 12699 18104 12708
rect 18052 12665 18061 12699
rect 18061 12665 18095 12699
rect 18095 12665 18104 12699
rect 18052 12656 18104 12665
rect 18512 12724 18564 12776
rect 19064 12724 19116 12776
rect 19432 12767 19484 12776
rect 19432 12733 19441 12767
rect 19441 12733 19475 12767
rect 19475 12733 19484 12767
rect 19432 12724 19484 12733
rect 19708 12767 19760 12776
rect 19708 12733 19742 12767
rect 19742 12733 19760 12767
rect 19708 12724 19760 12733
rect 20720 12724 20772 12776
rect 19340 12656 19392 12708
rect 20996 12656 21048 12708
rect 10784 12588 10836 12640
rect 10968 12631 11020 12640
rect 10968 12597 10977 12631
rect 10977 12597 11011 12631
rect 11011 12597 11020 12631
rect 10968 12588 11020 12597
rect 12256 12631 12308 12640
rect 12256 12597 12265 12631
rect 12265 12597 12299 12631
rect 12299 12597 12308 12631
rect 12256 12588 12308 12597
rect 14924 12631 14976 12640
rect 14924 12597 14933 12631
rect 14933 12597 14967 12631
rect 14967 12597 14976 12631
rect 14924 12588 14976 12597
rect 17960 12588 18012 12640
rect 19156 12588 19208 12640
rect 20812 12588 20864 12640
rect 21824 12792 21876 12844
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 22100 12656 22152 12708
rect 4322 12486 4374 12538
rect 4386 12486 4438 12538
rect 4450 12486 4502 12538
rect 4514 12486 4566 12538
rect 4578 12486 4630 12538
rect 5264 12384 5316 12436
rect 6460 12427 6512 12436
rect 6460 12393 6469 12427
rect 6469 12393 6503 12427
rect 6503 12393 6512 12427
rect 6460 12384 6512 12393
rect 6644 12384 6696 12436
rect 11428 12384 11480 12436
rect 11980 12384 12032 12436
rect 14004 12384 14056 12436
rect 14648 12384 14700 12436
rect 4896 12316 4948 12368
rect 7380 12316 7432 12368
rect 7932 12316 7984 12368
rect 8392 12359 8444 12368
rect 8392 12325 8401 12359
rect 8401 12325 8435 12359
rect 8435 12325 8444 12359
rect 8392 12316 8444 12325
rect 4252 12291 4304 12300
rect 4252 12257 4261 12291
rect 4261 12257 4295 12291
rect 4295 12257 4304 12291
rect 4252 12248 4304 12257
rect 8208 12291 8260 12300
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 8484 12291 8536 12300
rect 8484 12257 8493 12291
rect 8493 12257 8527 12291
rect 8527 12257 8536 12291
rect 8484 12248 8536 12257
rect 8576 12291 8628 12300
rect 8576 12257 8585 12291
rect 8585 12257 8619 12291
rect 8619 12257 8628 12291
rect 8576 12248 8628 12257
rect 9220 12291 9272 12300
rect 9220 12257 9229 12291
rect 9229 12257 9263 12291
rect 9263 12257 9272 12291
rect 9220 12248 9272 12257
rect 9772 12291 9824 12300
rect 9772 12257 9781 12291
rect 9781 12257 9815 12291
rect 9815 12257 9824 12291
rect 9772 12248 9824 12257
rect 12256 12316 12308 12368
rect 11520 12291 11572 12300
rect 11520 12257 11526 12291
rect 11526 12257 11560 12291
rect 11560 12257 11572 12291
rect 11520 12248 11572 12257
rect 16212 12316 16264 12368
rect 17316 12316 17368 12368
rect 17776 12316 17828 12368
rect 17960 12359 18012 12368
rect 17960 12325 17994 12359
rect 17994 12325 18012 12359
rect 17960 12316 18012 12325
rect 18052 12316 18104 12368
rect 19064 12427 19116 12436
rect 19064 12393 19073 12427
rect 19073 12393 19107 12427
rect 19107 12393 19116 12427
rect 19064 12384 19116 12393
rect 19156 12384 19208 12436
rect 20996 12427 21048 12436
rect 20996 12393 21005 12427
rect 21005 12393 21039 12427
rect 21039 12393 21048 12427
rect 20996 12384 21048 12393
rect 21640 12427 21692 12436
rect 21640 12393 21649 12427
rect 21649 12393 21683 12427
rect 21683 12393 21692 12427
rect 21640 12384 21692 12393
rect 20628 12316 20680 12368
rect 21364 12359 21416 12368
rect 21364 12325 21373 12359
rect 21373 12325 21407 12359
rect 21407 12325 21416 12359
rect 21364 12316 21416 12325
rect 22284 12316 22336 12368
rect 6828 12112 6880 12164
rect 9036 12180 9088 12232
rect 9680 12223 9732 12232
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 10692 12180 10744 12232
rect 14924 12248 14976 12300
rect 15108 12291 15160 12300
rect 15108 12257 15117 12291
rect 15117 12257 15151 12291
rect 15151 12257 15160 12291
rect 15108 12248 15160 12257
rect 16304 12291 16356 12300
rect 16304 12257 16313 12291
rect 16313 12257 16347 12291
rect 16347 12257 16356 12291
rect 16304 12248 16356 12257
rect 16948 12291 17000 12300
rect 16948 12257 16957 12291
rect 16957 12257 16991 12291
rect 16991 12257 17000 12291
rect 16948 12248 17000 12257
rect 20260 12248 20312 12300
rect 22008 12248 22060 12300
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 14556 12180 14608 12232
rect 16396 12223 16448 12232
rect 16396 12189 16405 12223
rect 16405 12189 16439 12223
rect 16439 12189 16448 12223
rect 16396 12180 16448 12189
rect 10876 12112 10928 12164
rect 8668 12044 8720 12096
rect 8944 12087 8996 12096
rect 8944 12053 8953 12087
rect 8953 12053 8987 12087
rect 8987 12053 8996 12087
rect 8944 12044 8996 12053
rect 14648 12044 14700 12096
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 18696 12180 18748 12232
rect 20444 12180 20496 12232
rect 19432 12044 19484 12096
rect 20168 12044 20220 12096
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 5632 11883 5684 11892
rect 5632 11849 5641 11883
rect 5641 11849 5675 11883
rect 5675 11849 5684 11883
rect 5632 11840 5684 11849
rect 8576 11840 8628 11892
rect 9588 11840 9640 11892
rect 11704 11840 11756 11892
rect 12072 11883 12124 11892
rect 12072 11849 12081 11883
rect 12081 11849 12115 11883
rect 12115 11849 12124 11883
rect 12072 11840 12124 11849
rect 14556 11840 14608 11892
rect 15108 11840 15160 11892
rect 17776 11840 17828 11892
rect 19800 11840 19852 11892
rect 21272 11883 21324 11892
rect 21272 11849 21281 11883
rect 21281 11849 21315 11883
rect 21315 11849 21324 11883
rect 21272 11840 21324 11849
rect 5540 11815 5592 11824
rect 5540 11781 5549 11815
rect 5549 11781 5583 11815
rect 5583 11781 5592 11815
rect 5540 11772 5592 11781
rect 19432 11772 19484 11824
rect 5264 11704 5316 11756
rect 6000 11704 6052 11756
rect 5172 11636 5224 11688
rect 8392 11679 8444 11688
rect 8392 11645 8401 11679
rect 8401 11645 8435 11679
rect 8435 11645 8444 11679
rect 8392 11636 8444 11645
rect 8668 11679 8720 11688
rect 8668 11645 8702 11679
rect 8702 11645 8720 11679
rect 8668 11636 8720 11645
rect 10692 11679 10744 11688
rect 10692 11645 10701 11679
rect 10701 11645 10735 11679
rect 10735 11645 10744 11679
rect 10692 11636 10744 11645
rect 10968 11679 11020 11688
rect 10968 11645 11002 11679
rect 11002 11645 11020 11679
rect 10968 11636 11020 11645
rect 14096 11636 14148 11688
rect 14280 11679 14332 11688
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 14648 11679 14700 11688
rect 14648 11645 14682 11679
rect 14682 11645 14700 11679
rect 13452 11568 13504 11620
rect 14648 11636 14700 11645
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 19156 11636 19208 11688
rect 20444 11636 20496 11688
rect 15016 11568 15068 11620
rect 18420 11568 18472 11620
rect 20260 11568 20312 11620
rect 20720 11636 20772 11688
rect 20996 11704 21048 11756
rect 21088 11636 21140 11688
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 19984 11500 20036 11552
rect 20720 11543 20772 11552
rect 20720 11509 20729 11543
rect 20729 11509 20763 11543
rect 20763 11509 20772 11543
rect 20720 11500 20772 11509
rect 20996 11500 21048 11552
rect 22284 11500 22336 11552
rect 22652 11500 22704 11552
rect 4322 11398 4374 11450
rect 4386 11398 4438 11450
rect 4450 11398 4502 11450
rect 4514 11398 4566 11450
rect 4578 11398 4630 11450
rect 5448 11296 5500 11348
rect 5172 11228 5224 11280
rect 5908 11271 5960 11280
rect 5908 11237 5917 11271
rect 5917 11237 5951 11271
rect 5951 11237 5960 11271
rect 5908 11228 5960 11237
rect 6276 11228 6328 11280
rect 8392 11296 8444 11348
rect 14280 11296 14332 11348
rect 5724 11092 5776 11144
rect 6000 11135 6052 11144
rect 6000 11101 6009 11135
rect 6009 11101 6043 11135
rect 6043 11101 6052 11135
rect 6000 11092 6052 11101
rect 10692 11228 10744 11280
rect 13820 11228 13872 11280
rect 8668 11160 8720 11212
rect 10968 11203 11020 11212
rect 10968 11169 10977 11203
rect 10977 11169 11011 11203
rect 11011 11169 11020 11203
rect 10968 11160 11020 11169
rect 11244 11203 11296 11212
rect 11244 11169 11278 11203
rect 11278 11169 11296 11203
rect 11244 11160 11296 11169
rect 13452 11203 13504 11212
rect 13452 11169 13461 11203
rect 13461 11169 13495 11203
rect 13495 11169 13504 11203
rect 13452 11160 13504 11169
rect 5632 11024 5684 11076
rect 7012 11024 7064 11076
rect 5724 10956 5776 11008
rect 9496 10999 9548 11008
rect 9496 10965 9505 10999
rect 9505 10965 9539 10999
rect 9539 10965 9548 10999
rect 9496 10956 9548 10965
rect 12348 10999 12400 11008
rect 12348 10965 12357 10999
rect 12357 10965 12391 10999
rect 12391 10965 12400 10999
rect 12348 10956 12400 10965
rect 14924 11296 14976 11348
rect 17316 11296 17368 11348
rect 20168 11296 20220 11348
rect 20812 11339 20864 11348
rect 20812 11305 20821 11339
rect 20821 11305 20855 11339
rect 20855 11305 20864 11339
rect 20812 11296 20864 11305
rect 21640 11296 21692 11348
rect 14924 11203 14976 11212
rect 14924 11169 14933 11203
rect 14933 11169 14967 11203
rect 14967 11169 14976 11203
rect 14924 11160 14976 11169
rect 15108 11203 15160 11212
rect 15108 11169 15117 11203
rect 15117 11169 15151 11203
rect 15151 11169 15160 11203
rect 15108 11160 15160 11169
rect 16212 11228 16264 11280
rect 17776 11228 17828 11280
rect 22008 11339 22060 11348
rect 22008 11305 22017 11339
rect 22017 11305 22051 11339
rect 22051 11305 22060 11339
rect 22008 11296 22060 11305
rect 22100 11296 22152 11348
rect 16580 11203 16632 11212
rect 16580 11169 16589 11203
rect 16589 11169 16623 11203
rect 16623 11169 16632 11203
rect 16580 11160 16632 11169
rect 16948 11160 17000 11212
rect 18420 11160 18472 11212
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 19708 11203 19760 11212
rect 19708 11169 19742 11203
rect 19742 11169 19760 11203
rect 19708 11160 19760 11169
rect 21732 11160 21784 11212
rect 16672 11135 16724 11144
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 20996 11092 21048 11144
rect 16396 11024 16448 11076
rect 16856 10999 16908 11008
rect 16856 10965 16865 10999
rect 16865 10965 16899 10999
rect 16899 10965 16908 10999
rect 16856 10956 16908 10965
rect 17040 10999 17092 11008
rect 17040 10965 17049 10999
rect 17049 10965 17083 10999
rect 17083 10965 17092 10999
rect 17040 10956 17092 10965
rect 20812 11024 20864 11076
rect 21364 11024 21416 11076
rect 17868 10999 17920 11008
rect 17868 10965 17877 10999
rect 17877 10965 17911 10999
rect 17911 10965 17920 10999
rect 17868 10956 17920 10965
rect 18236 10956 18288 11008
rect 21916 10956 21968 11008
rect 22008 10956 22060 11008
rect 22284 10999 22336 11008
rect 22284 10965 22293 10999
rect 22293 10965 22327 10999
rect 22327 10965 22336 10999
rect 22284 10956 22336 10965
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 5724 10752 5776 10804
rect 8668 10795 8720 10804
rect 8668 10761 8677 10795
rect 8677 10761 8711 10795
rect 8711 10761 8720 10795
rect 8668 10752 8720 10761
rect 9588 10795 9640 10804
rect 9588 10761 9597 10795
rect 9597 10761 9631 10795
rect 9631 10761 9640 10795
rect 9588 10752 9640 10761
rect 5172 10616 5224 10668
rect 5356 10616 5408 10668
rect 7196 10684 7248 10736
rect 11244 10752 11296 10804
rect 11428 10752 11480 10804
rect 12072 10795 12124 10804
rect 12072 10761 12081 10795
rect 12081 10761 12115 10795
rect 12115 10761 12124 10795
rect 12072 10752 12124 10761
rect 5908 10548 5960 10600
rect 6368 10591 6420 10600
rect 6368 10557 6377 10591
rect 6377 10557 6411 10591
rect 6411 10557 6420 10591
rect 6368 10548 6420 10557
rect 8944 10616 8996 10668
rect 9496 10616 9548 10668
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 10876 10659 10928 10668
rect 10876 10625 10885 10659
rect 10885 10625 10919 10659
rect 10919 10625 10928 10659
rect 10876 10616 10928 10625
rect 5080 10480 5132 10532
rect 5540 10480 5592 10532
rect 6092 10523 6144 10532
rect 6092 10489 6101 10523
rect 6101 10489 6135 10523
rect 6135 10489 6144 10523
rect 6092 10480 6144 10489
rect 7104 10523 7156 10532
rect 7104 10489 7113 10523
rect 7113 10489 7147 10523
rect 7147 10489 7156 10523
rect 7104 10480 7156 10489
rect 6276 10412 6328 10464
rect 8944 10480 8996 10532
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 7288 10412 7340 10421
rect 8852 10412 8904 10464
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 12440 10684 12492 10736
rect 11980 10591 12032 10600
rect 11980 10557 11989 10591
rect 11989 10557 12023 10591
rect 12023 10557 12032 10591
rect 11980 10548 12032 10557
rect 12072 10523 12124 10532
rect 12072 10489 12081 10523
rect 12081 10489 12115 10523
rect 12115 10489 12124 10523
rect 12348 10591 12400 10600
rect 12348 10557 12357 10591
rect 12357 10557 12391 10591
rect 12391 10557 12400 10591
rect 14280 10752 14332 10804
rect 17040 10752 17092 10804
rect 17224 10752 17276 10804
rect 19708 10752 19760 10804
rect 20720 10752 20772 10804
rect 20904 10752 20956 10804
rect 22560 10752 22612 10804
rect 22836 10795 22888 10804
rect 22836 10761 22845 10795
rect 22845 10761 22879 10795
rect 22879 10761 22888 10795
rect 22836 10752 22888 10761
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 21732 10684 21784 10736
rect 18696 10616 18748 10668
rect 12348 10548 12400 10557
rect 14832 10548 14884 10600
rect 15108 10591 15160 10600
rect 15108 10557 15117 10591
rect 15117 10557 15151 10591
rect 15151 10557 15160 10591
rect 15108 10548 15160 10557
rect 16212 10591 16264 10600
rect 16212 10557 16221 10591
rect 16221 10557 16255 10591
rect 16255 10557 16264 10591
rect 16212 10548 16264 10557
rect 16396 10548 16448 10600
rect 12072 10480 12124 10489
rect 16580 10523 16632 10532
rect 16580 10489 16589 10523
rect 16589 10489 16623 10523
rect 16623 10489 16632 10523
rect 16580 10480 16632 10489
rect 16856 10591 16908 10600
rect 16856 10557 16865 10591
rect 16865 10557 16899 10591
rect 16899 10557 16908 10591
rect 16856 10548 16908 10557
rect 18236 10591 18288 10600
rect 18236 10557 18254 10591
rect 18254 10557 18288 10591
rect 18236 10548 18288 10557
rect 23020 10591 23072 10600
rect 23020 10557 23029 10591
rect 23029 10557 23063 10591
rect 23063 10557 23072 10591
rect 23020 10548 23072 10557
rect 17776 10480 17828 10532
rect 19984 10523 20036 10532
rect 19984 10489 20011 10523
rect 20011 10489 20036 10523
rect 19984 10480 20036 10489
rect 20168 10523 20220 10532
rect 20168 10489 20177 10523
rect 20177 10489 20211 10523
rect 20211 10489 20220 10523
rect 20168 10480 20220 10489
rect 21088 10480 21140 10532
rect 21640 10480 21692 10532
rect 12440 10412 12492 10464
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 13636 10412 13688 10464
rect 14188 10412 14240 10464
rect 14740 10412 14792 10464
rect 16856 10412 16908 10464
rect 18972 10412 19024 10464
rect 22100 10412 22152 10464
rect 22468 10412 22520 10464
rect 4322 10310 4374 10362
rect 4386 10310 4438 10362
rect 4450 10310 4502 10362
rect 4514 10310 4566 10362
rect 4578 10310 4630 10362
rect 6368 10251 6420 10260
rect 6368 10217 6377 10251
rect 6377 10217 6411 10251
rect 6411 10217 6420 10251
rect 6368 10208 6420 10217
rect 7288 10251 7340 10260
rect 7288 10217 7313 10251
rect 7313 10217 7340 10251
rect 7288 10208 7340 10217
rect 3516 10140 3568 10192
rect 4160 10140 4212 10192
rect 5448 10140 5500 10192
rect 4988 10115 5040 10124
rect 4988 10081 4997 10115
rect 4997 10081 5031 10115
rect 5031 10081 5040 10115
rect 4988 10072 5040 10081
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 5264 10072 5316 10081
rect 5356 10115 5408 10124
rect 5356 10081 5365 10115
rect 5365 10081 5399 10115
rect 5399 10081 5408 10115
rect 5356 10072 5408 10081
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 6552 10072 6604 10124
rect 5632 10004 5684 10056
rect 7656 10115 7708 10124
rect 7656 10081 7665 10115
rect 7665 10081 7699 10115
rect 7699 10081 7708 10115
rect 7656 10072 7708 10081
rect 7932 10072 7984 10124
rect 8852 10208 8904 10260
rect 12348 10208 12400 10260
rect 17224 10208 17276 10260
rect 8484 10183 8536 10192
rect 8484 10149 8493 10183
rect 8493 10149 8527 10183
rect 8527 10149 8536 10183
rect 8484 10140 8536 10149
rect 9404 10183 9456 10192
rect 9404 10149 9413 10183
rect 9413 10149 9447 10183
rect 9447 10149 9456 10183
rect 9404 10140 9456 10149
rect 11520 10140 11572 10192
rect 17592 10251 17644 10260
rect 17592 10217 17601 10251
rect 17601 10217 17635 10251
rect 17635 10217 17644 10251
rect 17592 10208 17644 10217
rect 17868 10208 17920 10260
rect 22100 10208 22152 10260
rect 22192 10208 22244 10260
rect 8944 10115 8996 10124
rect 8116 10004 8168 10056
rect 4068 9936 4120 9988
rect 6368 9936 6420 9988
rect 3332 9868 3384 9920
rect 4252 9868 4304 9920
rect 6000 9868 6052 9920
rect 7012 9868 7064 9920
rect 7656 9936 7708 9988
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 11428 10115 11480 10124
rect 11428 10081 11437 10115
rect 11437 10081 11471 10115
rect 11471 10081 11480 10115
rect 11428 10072 11480 10081
rect 21088 10140 21140 10192
rect 22008 10140 22060 10192
rect 12072 10115 12124 10124
rect 12072 10081 12081 10115
rect 12081 10081 12115 10115
rect 12115 10081 12124 10115
rect 12072 10072 12124 10081
rect 8576 10004 8628 10056
rect 8852 10047 8904 10056
rect 8852 10013 8861 10047
rect 8861 10013 8895 10047
rect 8895 10013 8904 10047
rect 8852 10004 8904 10013
rect 12808 10072 12860 10124
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 14740 10115 14792 10124
rect 14740 10081 14749 10115
rect 14749 10081 14783 10115
rect 14783 10081 14792 10115
rect 14740 10072 14792 10081
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 16948 10072 17000 10124
rect 17408 10115 17460 10124
rect 17408 10081 17417 10115
rect 17417 10081 17451 10115
rect 17451 10081 17460 10115
rect 17408 10072 17460 10081
rect 17776 10115 17828 10124
rect 17776 10081 17785 10115
rect 17785 10081 17819 10115
rect 17819 10081 17828 10115
rect 17776 10072 17828 10081
rect 17868 10115 17920 10124
rect 17868 10081 17877 10115
rect 17877 10081 17911 10115
rect 17911 10081 17920 10115
rect 17868 10072 17920 10081
rect 20720 10115 20772 10124
rect 20720 10081 20729 10115
rect 20729 10081 20763 10115
rect 20763 10081 20772 10115
rect 20720 10072 20772 10081
rect 20904 10115 20956 10124
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 21180 10072 21232 10124
rect 21640 10115 21692 10124
rect 21640 10081 21649 10115
rect 21649 10081 21683 10115
rect 21683 10081 21692 10115
rect 21640 10072 21692 10081
rect 14188 10004 14240 10013
rect 21456 10047 21508 10056
rect 21456 10013 21465 10047
rect 21465 10013 21499 10047
rect 21499 10013 21508 10047
rect 21456 10004 21508 10013
rect 22744 10115 22796 10124
rect 22744 10081 22753 10115
rect 22753 10081 22787 10115
rect 22787 10081 22796 10115
rect 22744 10072 22796 10081
rect 7472 9911 7524 9920
rect 7472 9877 7481 9911
rect 7481 9877 7515 9911
rect 7515 9877 7524 9911
rect 7472 9868 7524 9877
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 8668 9868 8720 9920
rect 9128 9868 9180 9920
rect 14924 9936 14976 9988
rect 16672 9936 16724 9988
rect 17592 9936 17644 9988
rect 20812 9936 20864 9988
rect 22836 10004 22888 10056
rect 9312 9868 9364 9920
rect 11704 9911 11756 9920
rect 11704 9877 11713 9911
rect 11713 9877 11747 9911
rect 11747 9877 11756 9911
rect 11704 9868 11756 9877
rect 12348 9911 12400 9920
rect 12348 9877 12357 9911
rect 12357 9877 12391 9911
rect 12391 9877 12400 9911
rect 12348 9868 12400 9877
rect 14464 9868 14516 9920
rect 21272 9868 21324 9920
rect 21364 9868 21416 9920
rect 22376 9868 22428 9920
rect 22560 9911 22612 9920
rect 22560 9877 22569 9911
rect 22569 9877 22603 9911
rect 22603 9877 22612 9911
rect 22560 9868 22612 9877
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 3332 9707 3384 9716
rect 3332 9673 3341 9707
rect 3341 9673 3375 9707
rect 3375 9673 3384 9707
rect 3332 9664 3384 9673
rect 3516 9664 3568 9716
rect 4988 9664 5040 9716
rect 5448 9664 5500 9716
rect 6552 9707 6604 9716
rect 6552 9673 6561 9707
rect 6561 9673 6595 9707
rect 6595 9673 6604 9707
rect 6552 9664 6604 9673
rect 7840 9664 7892 9716
rect 8852 9664 8904 9716
rect 16672 9707 16724 9716
rect 16672 9673 16681 9707
rect 16681 9673 16715 9707
rect 16715 9673 16724 9707
rect 16672 9664 16724 9673
rect 20720 9707 20772 9716
rect 20720 9673 20729 9707
rect 20729 9673 20763 9707
rect 20763 9673 20772 9707
rect 20720 9664 20772 9673
rect 6368 9639 6420 9648
rect 6368 9605 6377 9639
rect 6377 9605 6411 9639
rect 6411 9605 6420 9639
rect 6368 9596 6420 9605
rect 8208 9639 8260 9648
rect 8208 9605 8217 9639
rect 8217 9605 8251 9639
rect 8251 9605 8260 9639
rect 8208 9596 8260 9605
rect 6092 9528 6144 9580
rect 8300 9528 8352 9580
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 4252 9503 4304 9512
rect 4252 9469 4286 9503
rect 4286 9469 4304 9503
rect 4252 9460 4304 9469
rect 5356 9460 5408 9512
rect 5540 9460 5592 9512
rect 6000 9392 6052 9444
rect 7196 9460 7248 9512
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 5264 9324 5316 9376
rect 5448 9324 5500 9376
rect 7656 9367 7708 9376
rect 7656 9333 7665 9367
rect 7665 9333 7699 9367
rect 7699 9333 7708 9367
rect 7656 9324 7708 9333
rect 8576 9460 8628 9512
rect 8944 9528 8996 9580
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 12348 9528 12400 9580
rect 13636 9571 13688 9580
rect 13636 9537 13645 9571
rect 13645 9537 13679 9571
rect 13679 9537 13688 9571
rect 13636 9528 13688 9537
rect 14464 9571 14516 9580
rect 14464 9537 14473 9571
rect 14473 9537 14507 9571
rect 14507 9537 14516 9571
rect 14464 9528 14516 9537
rect 14924 9571 14976 9580
rect 14924 9537 14933 9571
rect 14933 9537 14967 9571
rect 14967 9537 14976 9571
rect 14924 9528 14976 9537
rect 16580 9596 16632 9648
rect 21364 9664 21416 9716
rect 22836 9707 22888 9716
rect 22836 9673 22845 9707
rect 22845 9673 22879 9707
rect 22879 9673 22888 9707
rect 22836 9664 22888 9673
rect 9496 9460 9548 9512
rect 11336 9503 11388 9512
rect 11336 9469 11345 9503
rect 11345 9469 11379 9503
rect 11379 9469 11388 9503
rect 11336 9460 11388 9469
rect 13728 9503 13780 9512
rect 13728 9469 13737 9503
rect 13737 9469 13771 9503
rect 13771 9469 13780 9503
rect 13728 9460 13780 9469
rect 14372 9503 14424 9512
rect 14372 9469 14381 9503
rect 14381 9469 14415 9503
rect 14415 9469 14424 9503
rect 14372 9460 14424 9469
rect 15200 9460 15252 9512
rect 8484 9324 8536 9376
rect 8576 9324 8628 9376
rect 9404 9324 9456 9376
rect 11060 9324 11112 9376
rect 12256 9324 12308 9376
rect 16672 9460 16724 9512
rect 18052 9571 18104 9580
rect 18052 9537 18061 9571
rect 18061 9537 18095 9571
rect 18095 9537 18104 9571
rect 18052 9528 18104 9537
rect 18696 9528 18748 9580
rect 21180 9528 21232 9580
rect 17408 9460 17460 9512
rect 15476 9435 15528 9444
rect 15476 9401 15485 9435
rect 15485 9401 15519 9435
rect 15519 9401 15528 9435
rect 15476 9392 15528 9401
rect 16580 9367 16632 9376
rect 16580 9333 16589 9367
rect 16589 9333 16623 9367
rect 16623 9333 16632 9367
rect 16580 9324 16632 9333
rect 16764 9392 16816 9444
rect 19156 9435 19208 9444
rect 19156 9401 19165 9435
rect 19165 9401 19199 9435
rect 19199 9401 19208 9435
rect 19156 9392 19208 9401
rect 19616 9435 19668 9444
rect 19616 9401 19625 9435
rect 19625 9401 19659 9435
rect 19659 9401 19668 9435
rect 19616 9392 19668 9401
rect 21088 9460 21140 9512
rect 21364 9460 21416 9512
rect 21548 9460 21600 9512
rect 19892 9392 19944 9444
rect 20812 9392 20864 9444
rect 16856 9324 16908 9376
rect 18788 9367 18840 9376
rect 18788 9333 18797 9367
rect 18797 9333 18831 9367
rect 18831 9333 18840 9367
rect 18788 9324 18840 9333
rect 19524 9324 19576 9376
rect 21088 9324 21140 9376
rect 21824 9392 21876 9444
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 4988 9120 5040 9172
rect 4068 9052 4120 9104
rect 5080 9052 5132 9104
rect 7104 9052 7156 9104
rect 7656 9052 7708 9104
rect 15476 9120 15528 9172
rect 16764 9163 16816 9172
rect 16764 9129 16773 9163
rect 16773 9129 16807 9163
rect 16807 9129 16816 9163
rect 16764 9120 16816 9129
rect 17316 9120 17368 9172
rect 19892 9163 19944 9172
rect 19892 9129 19901 9163
rect 19901 9129 19935 9163
rect 19935 9129 19944 9163
rect 19892 9120 19944 9129
rect 15200 9052 15252 9104
rect 16488 9095 16540 9104
rect 16488 9061 16497 9095
rect 16497 9061 16531 9095
rect 16531 9061 16540 9095
rect 16488 9052 16540 9061
rect 16672 9052 16724 9104
rect 17408 9052 17460 9104
rect 17776 9095 17828 9104
rect 17776 9061 17785 9095
rect 17785 9061 17819 9095
rect 17819 9061 17828 9095
rect 17776 9052 17828 9061
rect 18788 9095 18840 9104
rect 18788 9061 18822 9095
rect 18822 9061 18840 9095
rect 18788 9052 18840 9061
rect 19432 9052 19484 9104
rect 20352 9120 20404 9172
rect 20904 9120 20956 9172
rect 21456 9120 21508 9172
rect 22560 9120 22612 9172
rect 5448 9027 5500 9036
rect 5448 8993 5457 9027
rect 5457 8993 5491 9027
rect 5491 8993 5500 9027
rect 5448 8984 5500 8993
rect 6092 9027 6144 9036
rect 6092 8993 6126 9027
rect 6126 8993 6144 9027
rect 5540 8916 5592 8968
rect 6092 8984 6144 8993
rect 7932 8984 7984 9036
rect 9128 8984 9180 9036
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 8300 8959 8352 8968
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 8300 8916 8352 8925
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 11704 8959 11756 8968
rect 11704 8925 11713 8959
rect 11713 8925 11747 8959
rect 11747 8925 11756 8959
rect 11704 8916 11756 8925
rect 3976 8780 4028 8832
rect 5632 8823 5684 8832
rect 5632 8789 5641 8823
rect 5641 8789 5675 8823
rect 5675 8789 5684 8823
rect 5632 8780 5684 8789
rect 14372 8984 14424 9036
rect 14556 8916 14608 8968
rect 18604 8984 18656 9036
rect 19708 8984 19760 9036
rect 20996 9052 21048 9104
rect 15016 8916 15068 8968
rect 16304 8959 16356 8968
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 18052 8916 18104 8968
rect 14464 8891 14516 8900
rect 14464 8857 14473 8891
rect 14473 8857 14507 8891
rect 14507 8857 14516 8891
rect 14464 8848 14516 8857
rect 16580 8848 16632 8900
rect 6828 8780 6880 8832
rect 8208 8780 8260 8832
rect 12256 8823 12308 8832
rect 12256 8789 12265 8823
rect 12265 8789 12299 8823
rect 12299 8789 12308 8823
rect 12256 8780 12308 8789
rect 16488 8780 16540 8832
rect 17868 8848 17920 8900
rect 20812 9027 20864 9036
rect 20812 8993 20821 9027
rect 20821 8993 20855 9027
rect 20855 8993 20864 9027
rect 20812 8984 20864 8993
rect 20076 8916 20128 8968
rect 21180 8984 21232 9036
rect 17592 8823 17644 8832
rect 17592 8789 17601 8823
rect 17601 8789 17635 8823
rect 17635 8789 17644 8823
rect 17592 8780 17644 8789
rect 20812 8780 20864 8832
rect 22008 8780 22060 8832
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 5632 8508 5684 8560
rect 6092 8619 6144 8628
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 10508 8576 10560 8628
rect 11336 8576 11388 8628
rect 13912 8619 13964 8628
rect 13912 8585 13921 8619
rect 13921 8585 13955 8619
rect 13955 8585 13964 8619
rect 13912 8576 13964 8585
rect 14372 8576 14424 8628
rect 17776 8619 17828 8628
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 20076 8619 20128 8628
rect 10876 8551 10928 8560
rect 10876 8517 10885 8551
rect 10885 8517 10919 8551
rect 10919 8517 10928 8551
rect 10876 8508 10928 8517
rect 10968 8508 11020 8560
rect 14648 8508 14700 8560
rect 15200 8508 15252 8560
rect 6368 8440 6420 8492
rect 7932 8415 7984 8424
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 8116 8372 8168 8381
rect 5080 8304 5132 8356
rect 7196 8304 7248 8356
rect 8484 8372 8536 8424
rect 9864 8440 9916 8492
rect 12992 8440 13044 8492
rect 10876 8372 10928 8424
rect 11520 8372 11572 8424
rect 11796 8372 11848 8424
rect 11888 8372 11940 8424
rect 14556 8440 14608 8492
rect 16304 8483 16356 8492
rect 16304 8449 16313 8483
rect 16313 8449 16347 8483
rect 16347 8449 16356 8483
rect 16304 8440 16356 8449
rect 17408 8440 17460 8492
rect 8392 8347 8444 8356
rect 8392 8313 8401 8347
rect 8401 8313 8435 8347
rect 8435 8313 8444 8347
rect 8392 8304 8444 8313
rect 8576 8347 8628 8356
rect 8576 8313 8585 8347
rect 8585 8313 8619 8347
rect 8619 8313 8628 8347
rect 8576 8304 8628 8313
rect 10692 8304 10744 8356
rect 11152 8304 11204 8356
rect 12348 8304 12400 8356
rect 13084 8304 13136 8356
rect 13728 8304 13780 8356
rect 14464 8304 14516 8356
rect 14556 8347 14608 8356
rect 14556 8313 14581 8347
rect 14581 8313 14608 8347
rect 14556 8304 14608 8313
rect 16488 8372 16540 8424
rect 17776 8372 17828 8424
rect 20076 8585 20085 8619
rect 20085 8585 20119 8619
rect 20119 8585 20128 8619
rect 20076 8576 20128 8585
rect 20904 8576 20956 8628
rect 21088 8576 21140 8628
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 19248 8372 19300 8424
rect 20812 8440 20864 8492
rect 15016 8304 15068 8356
rect 16948 8304 17000 8356
rect 4896 8236 4948 8288
rect 7564 8236 7616 8288
rect 7840 8236 7892 8288
rect 8852 8236 8904 8288
rect 8944 8279 8996 8288
rect 8944 8245 8953 8279
rect 8953 8245 8987 8279
rect 8987 8245 8996 8279
rect 8944 8236 8996 8245
rect 9772 8236 9824 8288
rect 10600 8236 10652 8288
rect 11060 8279 11112 8288
rect 11060 8245 11077 8279
rect 11077 8245 11112 8279
rect 11060 8236 11112 8245
rect 11612 8236 11664 8288
rect 11796 8279 11848 8288
rect 11796 8245 11805 8279
rect 11805 8245 11839 8279
rect 11839 8245 11848 8279
rect 11796 8236 11848 8245
rect 13176 8279 13228 8288
rect 13176 8245 13185 8279
rect 13185 8245 13219 8279
rect 13219 8245 13228 8279
rect 13176 8236 13228 8245
rect 13452 8236 13504 8288
rect 14280 8236 14332 8288
rect 14740 8279 14792 8288
rect 14740 8245 14749 8279
rect 14749 8245 14783 8279
rect 14783 8245 14792 8279
rect 14740 8236 14792 8245
rect 17960 8279 18012 8288
rect 17960 8245 17969 8279
rect 17969 8245 18003 8279
rect 18003 8245 18012 8279
rect 17960 8236 18012 8245
rect 18144 8279 18196 8288
rect 18144 8245 18153 8279
rect 18153 8245 18187 8279
rect 18187 8245 18196 8279
rect 18144 8236 18196 8245
rect 18788 8304 18840 8356
rect 19432 8304 19484 8356
rect 20996 8372 21048 8424
rect 21640 8372 21692 8424
rect 21916 8304 21968 8356
rect 20168 8279 20220 8288
rect 20168 8245 20177 8279
rect 20177 8245 20211 8279
rect 20211 8245 20220 8279
rect 20168 8236 20220 8245
rect 21088 8236 21140 8288
rect 21180 8279 21232 8288
rect 21180 8245 21189 8279
rect 21189 8245 21223 8279
rect 21223 8245 21232 8279
rect 21180 8236 21232 8245
rect 21272 8236 21324 8288
rect 21640 8236 21692 8288
rect 22652 8304 22704 8356
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 7196 8075 7248 8084
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 3516 7896 3568 7948
rect 5632 7964 5684 8016
rect 5724 7896 5776 7948
rect 7196 8041 7226 8075
rect 7226 8041 7248 8075
rect 7196 8032 7248 8041
rect 8392 8032 8444 8084
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 11336 8032 11388 8084
rect 11520 8075 11572 8084
rect 11520 8041 11529 8075
rect 11529 8041 11563 8075
rect 11563 8041 11572 8075
rect 11520 8032 11572 8041
rect 13084 8075 13136 8084
rect 13084 8041 13093 8075
rect 13093 8041 13127 8075
rect 13127 8041 13136 8075
rect 13084 8032 13136 8041
rect 13912 8032 13964 8084
rect 14280 8032 14332 8084
rect 7564 7964 7616 8016
rect 5448 7828 5500 7880
rect 7932 7964 7984 8016
rect 9956 7964 10008 8016
rect 10324 7964 10376 8016
rect 11704 7964 11756 8016
rect 12716 8007 12768 8016
rect 12716 7973 12725 8007
rect 12725 7973 12759 8007
rect 12759 7973 12768 8007
rect 12716 7964 12768 7973
rect 8024 7896 8076 7948
rect 8116 7939 8168 7948
rect 8116 7905 8125 7939
rect 8125 7905 8159 7939
rect 8159 7905 8168 7939
rect 8116 7896 8168 7905
rect 7196 7828 7248 7880
rect 10508 7939 10560 7948
rect 10508 7905 10517 7939
rect 10517 7905 10551 7939
rect 10551 7905 10560 7939
rect 10508 7896 10560 7905
rect 10600 7896 10652 7948
rect 8576 7828 8628 7880
rect 11060 7896 11112 7948
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 11612 7939 11664 7948
rect 11612 7905 11621 7939
rect 11621 7905 11655 7939
rect 11655 7905 11664 7939
rect 11612 7896 11664 7905
rect 12992 7939 13044 7948
rect 12992 7905 13001 7939
rect 13001 7905 13035 7939
rect 13035 7905 13044 7939
rect 12992 7896 13044 7905
rect 4068 7735 4120 7744
rect 4068 7701 4077 7735
rect 4077 7701 4111 7735
rect 4111 7701 4120 7735
rect 4068 7692 4120 7701
rect 4160 7692 4212 7744
rect 4896 7735 4948 7744
rect 4896 7701 4905 7735
rect 4905 7701 4939 7735
rect 4939 7701 4948 7735
rect 4896 7692 4948 7701
rect 5080 7735 5132 7744
rect 5080 7701 5089 7735
rect 5089 7701 5123 7735
rect 5123 7701 5132 7735
rect 5080 7692 5132 7701
rect 6552 7692 6604 7744
rect 7564 7760 7616 7812
rect 7932 7760 7984 7812
rect 9772 7760 9824 7812
rect 7840 7735 7892 7744
rect 7840 7701 7849 7735
rect 7849 7701 7883 7735
rect 7883 7701 7892 7735
rect 7840 7692 7892 7701
rect 8392 7692 8444 7744
rect 8760 7735 8812 7744
rect 8760 7701 8769 7735
rect 8769 7701 8803 7735
rect 8803 7701 8812 7735
rect 8760 7692 8812 7701
rect 8852 7692 8904 7744
rect 10232 7735 10284 7744
rect 10232 7701 10241 7735
rect 10241 7701 10275 7735
rect 10275 7701 10284 7735
rect 10232 7692 10284 7701
rect 10416 7692 10468 7744
rect 11152 7760 11204 7812
rect 14372 7896 14424 7948
rect 14648 8007 14700 8016
rect 14648 7973 14666 8007
rect 14666 7973 14700 8007
rect 15016 8075 15068 8084
rect 15016 8041 15025 8075
rect 15025 8041 15059 8075
rect 15059 8041 15068 8075
rect 15016 8032 15068 8041
rect 16672 8032 16724 8084
rect 14648 7964 14700 7973
rect 16488 8007 16540 8016
rect 16488 7973 16497 8007
rect 16497 7973 16531 8007
rect 16531 7973 16540 8007
rect 16488 7964 16540 7973
rect 18788 8075 18840 8084
rect 18788 8041 18797 8075
rect 18797 8041 18831 8075
rect 18831 8041 18840 8075
rect 18788 8032 18840 8041
rect 19524 8075 19576 8084
rect 19524 8041 19533 8075
rect 19533 8041 19567 8075
rect 19567 8041 19576 8075
rect 19524 8032 19576 8041
rect 19892 8032 19944 8084
rect 20812 8032 20864 8084
rect 21916 8032 21968 8084
rect 22652 8075 22704 8084
rect 22652 8041 22661 8075
rect 22661 8041 22695 8075
rect 22695 8041 22704 8075
rect 22652 8032 22704 8041
rect 18144 7964 18196 8016
rect 14924 7939 14976 7948
rect 14924 7905 14933 7939
rect 14933 7905 14967 7939
rect 14967 7905 14976 7939
rect 14924 7896 14976 7905
rect 17776 7896 17828 7948
rect 19524 7896 19576 7948
rect 20168 7964 20220 8016
rect 20996 7964 21048 8016
rect 21364 7964 21416 8016
rect 22008 7964 22060 8016
rect 21548 7939 21600 7948
rect 21548 7905 21582 7939
rect 21582 7905 21600 7939
rect 21548 7896 21600 7905
rect 21824 7896 21876 7948
rect 16488 7760 16540 7812
rect 16948 7803 17000 7812
rect 16948 7769 16957 7803
rect 16957 7769 16991 7803
rect 16991 7769 17000 7803
rect 16948 7760 17000 7769
rect 11796 7692 11848 7744
rect 12440 7735 12492 7744
rect 12440 7701 12449 7735
rect 12449 7701 12483 7735
rect 12483 7701 12492 7735
rect 12440 7692 12492 7701
rect 13360 7692 13412 7744
rect 14924 7692 14976 7744
rect 15384 7692 15436 7744
rect 17960 7692 18012 7744
rect 19156 7692 19208 7744
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 20720 7692 20772 7744
rect 22008 7692 22060 7744
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 3516 7531 3568 7540
rect 3516 7497 3525 7531
rect 3525 7497 3559 7531
rect 3559 7497 3568 7531
rect 3516 7488 3568 7497
rect 3608 7488 3660 7540
rect 4160 7488 4212 7540
rect 5632 7531 5684 7540
rect 5632 7497 5641 7531
rect 5641 7497 5675 7531
rect 5675 7497 5684 7531
rect 5632 7488 5684 7497
rect 6552 7531 6604 7540
rect 6552 7497 6561 7531
rect 6561 7497 6595 7531
rect 6595 7497 6604 7531
rect 6552 7488 6604 7497
rect 8116 7488 8168 7540
rect 8576 7488 8628 7540
rect 10232 7488 10284 7540
rect 11060 7488 11112 7540
rect 11244 7531 11296 7540
rect 11244 7497 11253 7531
rect 11253 7497 11287 7531
rect 11287 7497 11296 7531
rect 11244 7488 11296 7497
rect 11520 7488 11572 7540
rect 13176 7531 13228 7540
rect 13176 7497 13185 7531
rect 13185 7497 13219 7531
rect 13219 7497 13228 7531
rect 13176 7488 13228 7497
rect 13544 7488 13596 7540
rect 14464 7488 14516 7540
rect 15384 7531 15436 7540
rect 15384 7497 15393 7531
rect 15393 7497 15427 7531
rect 15427 7497 15436 7531
rect 15384 7488 15436 7497
rect 19524 7488 19576 7540
rect 21548 7488 21600 7540
rect 21824 7531 21876 7540
rect 21824 7497 21833 7531
rect 21833 7497 21867 7531
rect 21867 7497 21876 7531
rect 21824 7488 21876 7497
rect 4068 7420 4120 7472
rect 3332 7352 3384 7404
rect 3240 7284 3292 7336
rect 4068 7284 4120 7336
rect 4712 7216 4764 7268
rect 5724 7216 5776 7268
rect 5816 7259 5868 7268
rect 5816 7225 5825 7259
rect 5825 7225 5859 7259
rect 5859 7225 5868 7259
rect 5816 7216 5868 7225
rect 6000 7259 6052 7268
rect 6000 7225 6009 7259
rect 6009 7225 6043 7259
rect 6043 7225 6052 7259
rect 6000 7216 6052 7225
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 8944 7284 8996 7336
rect 12440 7327 12492 7336
rect 12440 7293 12458 7327
rect 12458 7293 12492 7327
rect 12440 7284 12492 7293
rect 3424 7148 3476 7200
rect 4160 7148 4212 7200
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 6552 7191 6604 7200
rect 6552 7157 6577 7191
rect 6577 7157 6604 7191
rect 8760 7216 8812 7268
rect 10232 7216 10284 7268
rect 10968 7216 11020 7268
rect 13452 7420 13504 7472
rect 6552 7148 6604 7157
rect 8024 7148 8076 7200
rect 11704 7148 11756 7200
rect 11888 7148 11940 7200
rect 13360 7284 13412 7336
rect 20076 7352 20128 7404
rect 13176 7191 13228 7200
rect 13176 7157 13201 7191
rect 13201 7157 13228 7191
rect 13176 7148 13228 7157
rect 14740 7284 14792 7336
rect 15200 7327 15252 7336
rect 15200 7293 15209 7327
rect 15209 7293 15243 7327
rect 15243 7293 15252 7327
rect 15200 7284 15252 7293
rect 19432 7327 19484 7336
rect 19432 7293 19441 7327
rect 19441 7293 19475 7327
rect 19475 7293 19484 7327
rect 19432 7284 19484 7293
rect 20904 7284 20956 7336
rect 21088 7284 21140 7336
rect 21640 7352 21692 7404
rect 21364 7327 21416 7336
rect 21364 7293 21373 7327
rect 21373 7293 21407 7327
rect 21407 7293 21416 7327
rect 21364 7284 21416 7293
rect 22744 7284 22796 7336
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 4252 6944 4304 6996
rect 3240 6876 3292 6928
rect 3792 6876 3844 6928
rect 3332 6808 3384 6860
rect 3240 6740 3292 6792
rect 3608 6672 3660 6724
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 4160 6808 4212 6860
rect 6552 6944 6604 6996
rect 7564 6987 7616 6996
rect 7564 6953 7573 6987
rect 7573 6953 7607 6987
rect 7607 6953 7616 6987
rect 7564 6944 7616 6953
rect 10232 6987 10284 6996
rect 10232 6953 10241 6987
rect 10241 6953 10275 6987
rect 10275 6953 10284 6987
rect 10232 6944 10284 6953
rect 12348 6987 12400 6996
rect 12348 6953 12357 6987
rect 12357 6953 12391 6987
rect 12391 6953 12400 6987
rect 12348 6944 12400 6953
rect 13176 6944 13228 6996
rect 5540 6876 5592 6928
rect 7196 6919 7248 6928
rect 7196 6885 7205 6919
rect 7205 6885 7239 6919
rect 7239 6885 7248 6919
rect 7196 6876 7248 6885
rect 7288 6876 7340 6928
rect 9956 6876 10008 6928
rect 13544 6919 13596 6928
rect 13544 6885 13553 6919
rect 13553 6885 13587 6919
rect 13587 6885 13596 6919
rect 13544 6876 13596 6885
rect 5816 6851 5868 6860
rect 5816 6817 5825 6851
rect 5825 6817 5859 6851
rect 5859 6817 5868 6851
rect 5816 6808 5868 6817
rect 6000 6851 6052 6860
rect 6000 6817 6009 6851
rect 6009 6817 6043 6851
rect 6043 6817 6052 6851
rect 6000 6808 6052 6817
rect 8392 6808 8444 6860
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 10876 6808 10928 6860
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 11060 6808 11112 6860
rect 12992 6808 13044 6860
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 5448 6740 5500 6792
rect 4160 6672 4212 6724
rect 5540 6604 5592 6656
rect 10416 6647 10468 6656
rect 10416 6613 10425 6647
rect 10425 6613 10459 6647
rect 10459 6613 10468 6647
rect 10416 6604 10468 6613
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 3424 6443 3476 6452
rect 3424 6409 3433 6443
rect 3433 6409 3467 6443
rect 3467 6409 3476 6443
rect 3424 6400 3476 6409
rect 4068 6400 4120 6452
rect 3240 6196 3292 6248
rect 4160 6196 4212 6248
rect 6000 6400 6052 6452
rect 10324 6400 10376 6452
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 6828 6264 6880 6316
rect 3332 6128 3384 6180
rect 5080 6196 5132 6248
rect 10692 6196 10744 6248
rect 11612 6128 11664 6180
rect 5816 6060 5868 6112
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 5816 5856 5868 5908
rect 3516 5788 3568 5840
rect 5724 5720 5776 5772
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 22744 4131 22796 4140
rect 22744 4097 22753 4131
rect 22753 4097 22787 4131
rect 22787 4097 22796 4131
rect 22744 4088 22796 4097
rect 22928 3995 22980 4004
rect 22928 3961 22937 3995
rect 22937 3961 22971 3995
rect 22971 3961 22980 3995
rect 22928 3952 22980 3961
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
<< metal2 >>
rect 1674 23746 1730 24000
rect 1674 23718 1808 23746
rect 1674 23600 1730 23718
rect 1780 23186 1808 23718
rect 4618 23610 4674 24000
rect 7562 23746 7618 24000
rect 7562 23718 7880 23746
rect 4618 23600 4752 23610
rect 7562 23600 7618 23718
rect 4632 23582 4752 23600
rect 4322 23420 4630 23429
rect 4322 23418 4328 23420
rect 4384 23418 4408 23420
rect 4464 23418 4488 23420
rect 4544 23418 4568 23420
rect 4624 23418 4630 23420
rect 4384 23366 4386 23418
rect 4566 23366 4568 23418
rect 4322 23364 4328 23366
rect 4384 23364 4408 23366
rect 4464 23364 4488 23366
rect 4544 23364 4568 23366
rect 4624 23364 4630 23366
rect 4322 23355 4630 23364
rect 4724 23254 4752 23582
rect 4712 23248 4764 23254
rect 4712 23190 4764 23196
rect 7852 23186 7880 23718
rect 10506 23600 10562 24000
rect 13450 23746 13506 24000
rect 16394 23746 16450 24000
rect 13450 23718 13584 23746
rect 13450 23600 13506 23718
rect 10520 23254 10548 23600
rect 10508 23248 10560 23254
rect 10508 23190 10560 23196
rect 13556 23186 13584 23718
rect 16394 23718 16528 23746
rect 16394 23600 16450 23718
rect 16500 23186 16528 23718
rect 19338 23600 19394 24000
rect 22282 23600 22338 24000
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 1768 23180 1820 23186
rect 1768 23122 1820 23128
rect 5356 23180 5408 23186
rect 5356 23122 5408 23128
rect 6460 23180 6512 23186
rect 6460 23122 6512 23128
rect 6920 23180 6972 23186
rect 6920 23122 6972 23128
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 8668 23180 8720 23186
rect 8668 23122 8720 23128
rect 8852 23180 8904 23186
rect 8852 23122 8904 23128
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 16488 23180 16540 23186
rect 16488 23122 16540 23128
rect 5368 22982 5396 23122
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 5356 22976 5408 22982
rect 5356 22918 5408 22924
rect 3662 22876 3970 22885
rect 3662 22874 3668 22876
rect 3724 22874 3748 22876
rect 3804 22874 3828 22876
rect 3884 22874 3908 22876
rect 3964 22874 3970 22876
rect 3724 22822 3726 22874
rect 3906 22822 3908 22874
rect 3662 22820 3668 22822
rect 3724 22820 3748 22822
rect 3804 22820 3828 22822
rect 3884 22820 3908 22822
rect 3964 22820 3970 22822
rect 3662 22811 3970 22820
rect 4908 22710 4936 22918
rect 4712 22704 4764 22710
rect 4712 22646 4764 22652
rect 4896 22704 4948 22710
rect 4896 22646 4948 22652
rect 4252 22500 4304 22506
rect 4252 22442 4304 22448
rect 4264 22166 4292 22442
rect 4322 22332 4630 22341
rect 4322 22330 4328 22332
rect 4384 22330 4408 22332
rect 4464 22330 4488 22332
rect 4544 22330 4568 22332
rect 4624 22330 4630 22332
rect 4384 22278 4386 22330
rect 4566 22278 4568 22330
rect 4322 22276 4328 22278
rect 4384 22276 4408 22278
rect 4464 22276 4488 22278
rect 4544 22276 4568 22278
rect 4624 22276 4630 22278
rect 4322 22267 4630 22276
rect 4252 22160 4304 22166
rect 4252 22102 4304 22108
rect 3662 21788 3970 21797
rect 3662 21786 3668 21788
rect 3724 21786 3748 21788
rect 3804 21786 3828 21788
rect 3884 21786 3908 21788
rect 3964 21786 3970 21788
rect 3724 21734 3726 21786
rect 3906 21734 3908 21786
rect 3662 21732 3668 21734
rect 3724 21732 3748 21734
rect 3804 21732 3828 21734
rect 3884 21732 3908 21734
rect 3964 21732 3970 21734
rect 3662 21723 3970 21732
rect 3662 20700 3970 20709
rect 3662 20698 3668 20700
rect 3724 20698 3748 20700
rect 3804 20698 3828 20700
rect 3884 20698 3908 20700
rect 3964 20698 3970 20700
rect 3724 20646 3726 20698
rect 3906 20646 3908 20698
rect 3662 20644 3668 20646
rect 3724 20644 3748 20646
rect 3804 20644 3828 20646
rect 3884 20644 3908 20646
rect 3964 20644 3970 20646
rect 3662 20635 3970 20644
rect 4264 20398 4292 22102
rect 4724 21962 4752 22646
rect 5368 22574 5396 22918
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 5356 22568 5408 22574
rect 5356 22510 5408 22516
rect 5908 22568 5960 22574
rect 5908 22510 5960 22516
rect 6368 22568 6420 22574
rect 6368 22510 6420 22516
rect 4816 22234 4844 22510
rect 4804 22228 4856 22234
rect 4804 22170 4856 22176
rect 4816 22094 4844 22170
rect 5632 22160 5684 22166
rect 5632 22102 5684 22108
rect 4816 22066 4936 22094
rect 4712 21956 4764 21962
rect 4712 21898 4764 21904
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4322 21244 4630 21253
rect 4322 21242 4328 21244
rect 4384 21242 4408 21244
rect 4464 21242 4488 21244
rect 4544 21242 4568 21244
rect 4624 21242 4630 21244
rect 4384 21190 4386 21242
rect 4566 21190 4568 21242
rect 4322 21188 4328 21190
rect 4384 21188 4408 21190
rect 4464 21188 4488 21190
rect 4544 21188 4568 21190
rect 4624 21188 4630 21190
rect 4322 21179 4630 21188
rect 4724 21010 4752 21286
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 4620 20392 4672 20398
rect 4724 20380 4752 20946
rect 4672 20352 4752 20380
rect 4620 20334 4672 20340
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 3662 19612 3970 19621
rect 3662 19610 3668 19612
rect 3724 19610 3748 19612
rect 3804 19610 3828 19612
rect 3884 19610 3908 19612
rect 3964 19610 3970 19612
rect 3724 19558 3726 19610
rect 3906 19558 3908 19610
rect 3662 19556 3668 19558
rect 3724 19556 3748 19558
rect 3804 19556 3828 19558
rect 3884 19556 3908 19558
rect 3964 19556 3970 19558
rect 3662 19547 3970 19556
rect 4172 19378 4200 19926
rect 4264 19718 4292 20198
rect 4322 20156 4630 20165
rect 4322 20154 4328 20156
rect 4384 20154 4408 20156
rect 4464 20154 4488 20156
rect 4544 20154 4568 20156
rect 4624 20154 4630 20156
rect 4384 20102 4386 20154
rect 4566 20102 4568 20154
rect 4322 20100 4328 20102
rect 4384 20100 4408 20102
rect 4464 20100 4488 20102
rect 4544 20100 4568 20102
rect 4624 20100 4630 20102
rect 4322 20091 4630 20100
rect 4344 19780 4396 19786
rect 4344 19722 4396 19728
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4264 19310 4292 19654
rect 4356 19310 4384 19722
rect 4724 19378 4752 20352
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 4816 19718 4844 20334
rect 4908 19990 4936 22066
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 4896 19984 4948 19990
rect 4896 19926 4948 19932
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4816 19514 4844 19654
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 4344 19304 4396 19310
rect 4804 19304 4856 19310
rect 4344 19246 4396 19252
rect 4802 19272 4804 19281
rect 4856 19272 4858 19281
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 3662 18459 3970 18468
rect 4264 18306 4292 19246
rect 4802 19207 4858 19216
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4322 19068 4630 19077
rect 4322 19066 4328 19068
rect 4384 19066 4408 19068
rect 4464 19066 4488 19068
rect 4544 19066 4568 19068
rect 4624 19066 4630 19068
rect 4384 19014 4386 19066
rect 4566 19014 4568 19066
rect 4322 19012 4328 19014
rect 4384 19012 4408 19014
rect 4464 19012 4488 19014
rect 4544 19012 4568 19014
rect 4624 19012 4630 19014
rect 4322 19003 4630 19012
rect 4160 18284 4212 18290
rect 4264 18278 4384 18306
rect 4160 18226 4212 18232
rect 4172 17882 4200 18226
rect 4356 18154 4384 18278
rect 4620 18216 4672 18222
rect 4672 18164 4752 18170
rect 4620 18158 4752 18164
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4344 18148 4396 18154
rect 4632 18142 4752 18158
rect 4344 18090 4396 18096
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 4080 15570 4108 16662
rect 4172 16658 4200 17818
rect 4264 17338 4292 18090
rect 4322 17980 4630 17989
rect 4322 17978 4328 17980
rect 4384 17978 4408 17980
rect 4464 17978 4488 17980
rect 4544 17978 4568 17980
rect 4624 17978 4630 17980
rect 4384 17926 4386 17978
rect 4566 17926 4568 17978
rect 4322 17924 4328 17926
rect 4384 17924 4408 17926
rect 4464 17924 4488 17926
rect 4544 17924 4568 17926
rect 4624 17924 4630 17926
rect 4322 17915 4630 17924
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4264 16794 4292 17274
rect 4356 17066 4384 17682
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4448 17134 4476 17614
rect 4632 17218 4660 17682
rect 4724 17542 4752 18142
rect 4816 17814 4844 19110
rect 4908 18222 4936 19926
rect 5000 19242 5028 21966
rect 5448 21888 5500 21894
rect 5448 21830 5500 21836
rect 5460 21690 5488 21830
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 5092 20058 5120 20334
rect 5172 20324 5224 20330
rect 5172 20266 5224 20272
rect 5080 20052 5132 20058
rect 5080 19994 5132 20000
rect 5184 19922 5212 20266
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 5184 19514 5212 19858
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5172 19372 5224 19378
rect 5224 19332 5304 19360
rect 5172 19314 5224 19320
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5184 18358 5212 18770
rect 5172 18352 5224 18358
rect 5172 18294 5224 18300
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4804 17808 4856 17814
rect 4804 17750 4856 17756
rect 4908 17678 4936 18158
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4724 17338 4752 17478
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4632 17190 4752 17218
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 4448 16998 4476 17070
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4322 16892 4630 16901
rect 4322 16890 4328 16892
rect 4384 16890 4408 16892
rect 4464 16890 4488 16892
rect 4544 16890 4568 16892
rect 4624 16890 4630 16892
rect 4384 16838 4386 16890
rect 4566 16838 4568 16890
rect 4322 16836 4328 16838
rect 4384 16836 4408 16838
rect 4464 16836 4488 16838
rect 4544 16836 4568 16838
rect 4624 16836 4630 16838
rect 4322 16827 4630 16836
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4724 16726 4752 17190
rect 5000 17134 5028 18226
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 5092 17066 5120 18090
rect 5080 17060 5132 17066
rect 5080 17002 5132 17008
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4264 15706 4292 16526
rect 4322 15804 4630 15813
rect 4322 15802 4328 15804
rect 4384 15802 4408 15804
rect 4464 15802 4488 15804
rect 4544 15802 4568 15804
rect 4624 15802 4630 15804
rect 4384 15750 4386 15802
rect 4566 15750 4568 15802
rect 4322 15748 4328 15750
rect 4384 15748 4408 15750
rect 4464 15748 4488 15750
rect 4544 15748 4568 15750
rect 4624 15748 4630 15750
rect 4322 15739 4630 15748
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4080 15450 4108 15506
rect 4724 15502 4752 16526
rect 5092 16522 5120 17002
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 16658 5212 16934
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 5080 16516 5132 16522
rect 5080 16458 5132 16464
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4712 15496 4764 15502
rect 4080 15422 4200 15450
rect 4712 15438 4764 15444
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 4172 15162 4200 15422
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4816 14958 4844 15642
rect 5092 15570 5120 16458
rect 5276 16046 5304 19332
rect 5460 19310 5488 21626
rect 5644 21010 5672 22102
rect 5920 21078 5948 22510
rect 6276 21480 6328 21486
rect 6380 21468 6408 22510
rect 6472 22166 6500 23122
rect 6932 22778 6960 23122
rect 7472 23112 7524 23118
rect 7472 23054 7524 23060
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 7484 22574 7512 23054
rect 8116 23044 8168 23050
rect 8116 22986 8168 22992
rect 7472 22568 7524 22574
rect 7472 22510 7524 22516
rect 7564 22568 7616 22574
rect 7564 22510 7616 22516
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 7196 22500 7248 22506
rect 7196 22442 7248 22448
rect 6460 22160 6512 22166
rect 6460 22102 6512 22108
rect 6736 22160 6788 22166
rect 6736 22102 6788 22108
rect 6748 21486 6776 22102
rect 7208 22098 7236 22442
rect 7576 22438 7604 22510
rect 7564 22432 7616 22438
rect 7564 22374 7616 22380
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 7196 22092 7248 22098
rect 7576 22094 7604 22374
rect 7196 22034 7248 22040
rect 7484 22066 7604 22094
rect 6840 21622 6868 22034
rect 7484 21962 7512 22066
rect 6920 21956 6972 21962
rect 6920 21898 6972 21904
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 6828 21616 6880 21622
rect 6828 21558 6880 21564
rect 6840 21486 6868 21558
rect 6328 21440 6408 21468
rect 6276 21422 6328 21428
rect 5908 21072 5960 21078
rect 5908 21014 5960 21020
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5644 20398 5672 20946
rect 6380 20942 6408 21440
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 6828 21480 6880 21486
rect 6828 21422 6880 21428
rect 6748 21146 6776 21422
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6368 20936 6420 20942
rect 6090 20904 6146 20913
rect 6368 20878 6420 20884
rect 6090 20839 6146 20848
rect 6736 20868 6788 20874
rect 6104 20806 6132 20839
rect 6736 20810 6788 20816
rect 6092 20800 6144 20806
rect 6092 20742 6144 20748
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6104 20398 6132 20742
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 6012 19922 6040 20198
rect 6000 19916 6052 19922
rect 6000 19858 6052 19864
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5448 19304 5500 19310
rect 5552 19281 5580 19654
rect 6012 19310 6040 19858
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6000 19304 6052 19310
rect 5448 19246 5500 19252
rect 5538 19272 5594 19281
rect 5460 18834 5488 19246
rect 6000 19246 6052 19252
rect 6104 19242 6132 19790
rect 5538 19207 5594 19216
rect 6092 19236 6144 19242
rect 6092 19178 6144 19184
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5644 18222 5672 18838
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5644 17814 5672 18158
rect 5632 17808 5684 17814
rect 5552 17756 5632 17762
rect 5552 17750 5684 17756
rect 5552 17734 5672 17750
rect 5552 17202 5580 17734
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5644 17338 5672 17614
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5552 16810 5580 17138
rect 5460 16794 5580 16810
rect 5448 16788 5580 16794
rect 5500 16782 5580 16788
rect 5448 16730 5500 16736
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5368 16114 5396 16390
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5828 15570 5856 18770
rect 5920 17746 5948 19110
rect 6104 18698 6132 19178
rect 6092 18692 6144 18698
rect 6092 18634 6144 18640
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 6012 17202 6040 18022
rect 6104 17610 6132 18158
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6092 17604 6144 17610
rect 6092 17546 6144 17552
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6104 17134 6132 17546
rect 6288 17202 6316 18022
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5092 15450 5120 15506
rect 5092 15422 5212 15450
rect 6012 15434 6040 15506
rect 6104 15502 6132 17070
rect 6288 16658 6316 17138
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 5184 14958 5212 15422
rect 6000 15428 6052 15434
rect 6000 15370 6052 15376
rect 6012 15094 6040 15370
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 6104 15026 6132 15438
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4264 14550 4292 14758
rect 4322 14716 4630 14725
rect 4322 14714 4328 14716
rect 4384 14714 4408 14716
rect 4464 14714 4488 14716
rect 4544 14714 4568 14716
rect 4624 14714 4630 14716
rect 4384 14662 4386 14714
rect 4566 14662 4568 14714
rect 4322 14660 4328 14662
rect 4384 14660 4408 14662
rect 4464 14660 4488 14662
rect 4544 14660 4568 14662
rect 4624 14660 4630 14662
rect 4322 14651 4630 14660
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 4322 13628 4630 13637
rect 4322 13626 4328 13628
rect 4384 13626 4408 13628
rect 4464 13626 4488 13628
rect 4544 13626 4568 13628
rect 4624 13626 4630 13628
rect 4384 13574 4386 13626
rect 4566 13574 4568 13626
rect 4322 13572 4328 13574
rect 4384 13572 4408 13574
rect 4464 13572 4488 13574
rect 4544 13572 4568 13574
rect 4624 13572 4630 13574
rect 4322 13563 4630 13572
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4264 12306 4292 12650
rect 4322 12540 4630 12549
rect 4322 12538 4328 12540
rect 4384 12538 4408 12540
rect 4464 12538 4488 12540
rect 4544 12538 4568 12540
rect 4624 12538 4630 12540
rect 4384 12486 4386 12538
rect 4566 12486 4568 12538
rect 4322 12484 4328 12486
rect 4384 12484 4408 12486
rect 4464 12484 4488 12486
rect 4544 12484 4568 12486
rect 4624 12484 4630 12486
rect 4322 12475 4630 12484
rect 4908 12374 4936 13126
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 5184 11694 5212 14010
rect 5460 13802 5488 14894
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 14278 5672 14758
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5354 13696 5410 13705
rect 5354 13631 5410 13640
rect 5368 13530 5396 13631
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5276 12442 5304 13330
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5276 11762 5304 12378
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 4322 11452 4630 11461
rect 4322 11450 4328 11452
rect 4384 11450 4408 11452
rect 4464 11450 4488 11452
rect 4544 11450 4568 11452
rect 4624 11450 4630 11452
rect 4384 11398 4386 11450
rect 4566 11398 4568 11450
rect 4322 11396 4328 11398
rect 4384 11396 4408 11398
rect 4464 11396 4488 11398
rect 4544 11396 4568 11398
rect 4624 11396 4630 11398
rect 4322 11387 4630 11396
rect 5184 11286 5212 11630
rect 5460 11354 5488 12650
rect 5644 11898 5672 14214
rect 6380 13530 6408 20742
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6564 18426 6592 18702
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5828 12782 5856 13126
rect 6196 12986 6224 13330
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 5184 10674 5212 11222
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 4322 10364 4630 10373
rect 4322 10362 4328 10364
rect 4384 10362 4408 10364
rect 4464 10362 4488 10364
rect 4544 10362 4568 10364
rect 4624 10362 4630 10364
rect 4384 10310 4386 10362
rect 4566 10310 4568 10362
rect 4322 10308 4328 10310
rect 4384 10308 4408 10310
rect 4464 10308 4488 10310
rect 4544 10308 4568 10310
rect 4624 10308 4630 10310
rect 4322 10299 4630 10308
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3344 9722 3372 9862
rect 3528 9722 3556 10134
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3988 8838 4016 9454
rect 4080 9110 4108 9930
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3528 7546 3556 7890
rect 4172 7750 4200 10134
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4264 9518 4292 9862
rect 5000 9722 5028 10066
rect 4988 9716 5040 9722
rect 4988 9658 5040 9664
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 5000 9178 5028 9658
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5092 9110 5120 10474
rect 5368 10130 5396 10610
rect 5552 10538 5580 11766
rect 5644 11234 5672 11834
rect 5920 11286 5948 12922
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6472 12442 6500 12650
rect 6656 12442 6684 20742
rect 6748 20398 6776 20810
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6840 18902 6868 21286
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6840 18766 6868 18838
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6932 18698 6960 21898
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7668 21486 7696 21626
rect 8036 21486 8064 22510
rect 8128 22098 8156 22986
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 8220 22642 8248 22714
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8116 21956 8168 21962
rect 8116 21898 8168 21904
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 7380 21412 7432 21418
rect 7380 21354 7432 21360
rect 7392 21010 7420 21354
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7024 20602 7052 20878
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 7668 20534 7696 21422
rect 8036 21146 8064 21422
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8128 20942 8156 21898
rect 8220 21622 8248 22578
rect 8312 22506 8340 23054
rect 8680 22778 8708 23122
rect 8668 22772 8720 22778
rect 8668 22714 8720 22720
rect 8484 22704 8536 22710
rect 8484 22646 8536 22652
rect 8300 22500 8352 22506
rect 8300 22442 8352 22448
rect 8496 22094 8524 22646
rect 8576 22432 8628 22438
rect 8680 22420 8708 22714
rect 8864 22574 8892 23122
rect 9220 23112 9272 23118
rect 9220 23054 9272 23060
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 9036 23044 9088 23050
rect 9036 22986 9088 22992
rect 9048 22710 9076 22986
rect 9036 22704 9088 22710
rect 9036 22646 9088 22652
rect 8760 22568 8812 22574
rect 8760 22510 8812 22516
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8628 22392 8708 22420
rect 8576 22374 8628 22380
rect 8496 22066 8616 22094
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8208 21616 8260 21622
rect 8208 21558 8260 21564
rect 8312 21486 8340 21966
rect 8588 21486 8616 22066
rect 8680 21486 8708 22392
rect 8772 21690 8800 22510
rect 8944 22432 8996 22438
rect 8944 22374 8996 22380
rect 8956 22234 8984 22374
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 8852 22024 8904 22030
rect 8852 21966 8904 21972
rect 8864 21894 8892 21966
rect 8852 21888 8904 21894
rect 8852 21830 8904 21836
rect 8760 21684 8812 21690
rect 8760 21626 8812 21632
rect 8956 21486 8984 22170
rect 9048 22166 9076 22646
rect 9036 22160 9088 22166
rect 9036 22102 9088 22108
rect 8300 21480 8352 21486
rect 8300 21422 8352 21428
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8312 21010 8340 21422
rect 8588 21010 8616 21422
rect 8758 21040 8814 21049
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8576 21004 8628 21010
rect 8758 20975 8814 20984
rect 8576 20946 8628 20952
rect 8116 20936 8168 20942
rect 8116 20878 8168 20884
rect 8772 20874 8800 20975
rect 8760 20868 8812 20874
rect 8760 20810 8812 20816
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 7656 20528 7708 20534
rect 7656 20470 7708 20476
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 7024 19310 7052 19858
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 7116 19378 7144 19722
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7472 19304 7524 19310
rect 7472 19246 7524 19252
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 7208 18630 7236 19246
rect 7484 18970 7512 19246
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7208 18154 7236 18566
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 7196 18148 7248 18154
rect 7196 18090 7248 18096
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6748 15502 6776 16050
rect 7024 16046 7052 18090
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 7392 17134 7420 17682
rect 7484 17270 7512 17682
rect 7472 17264 7524 17270
rect 7472 17206 7524 17212
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7576 16658 7604 19790
rect 7852 19310 7880 20742
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 7944 18970 7972 19178
rect 8036 18970 8064 19246
rect 7932 18964 7984 18970
rect 7932 18906 7984 18912
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8116 18692 8168 18698
rect 8116 18634 8168 18640
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6932 15162 6960 15914
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 7024 14958 7052 15370
rect 7116 15026 7144 16118
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7208 15502 7236 15982
rect 7576 15570 7604 16594
rect 8024 15972 8076 15978
rect 8024 15914 8076 15920
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6932 13938 6960 14758
rect 7208 14482 7236 15098
rect 8036 14550 8064 15914
rect 8024 14544 8076 14550
rect 8024 14486 8076 14492
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 7208 13870 7236 14418
rect 8128 14414 8156 18634
rect 8312 14482 8340 20742
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8772 18902 8800 19246
rect 8760 18896 8812 18902
rect 8760 18838 8812 18844
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8496 18154 8524 18770
rect 8772 18358 8800 18838
rect 9048 18834 9076 22102
rect 9232 21486 9260 23054
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9324 22574 9352 22714
rect 9508 22574 9536 23054
rect 9312 22568 9364 22574
rect 9312 22510 9364 22516
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 9324 21894 9352 22374
rect 9600 22234 9628 22510
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9876 22098 9904 22442
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9232 21078 9260 21422
rect 9220 21072 9272 21078
rect 9220 21014 9272 21020
rect 9220 20936 9272 20942
rect 9220 20878 9272 20884
rect 9232 20806 9260 20878
rect 9220 20800 9272 20806
rect 9220 20742 9272 20748
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 9048 18358 9076 18770
rect 8760 18352 8812 18358
rect 8760 18294 8812 18300
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 9324 18222 9352 21830
rect 9416 20874 9444 21966
rect 9770 21584 9826 21593
rect 9770 21519 9826 21528
rect 9496 21480 9548 21486
rect 9496 21422 9548 21428
rect 9508 21162 9536 21422
rect 9508 21146 9628 21162
rect 9508 21140 9640 21146
rect 9508 21134 9588 21140
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9508 18154 9536 21134
rect 9588 21082 9640 21088
rect 9784 21078 9812 21519
rect 10152 21486 10180 23054
rect 11336 22976 11388 22982
rect 11336 22918 11388 22924
rect 14924 22976 14976 22982
rect 14924 22918 14976 22924
rect 10600 22568 10652 22574
rect 10600 22510 10652 22516
rect 10506 21992 10562 22001
rect 10506 21927 10562 21936
rect 10322 21584 10378 21593
rect 10322 21519 10378 21528
rect 10336 21486 10364 21519
rect 10140 21480 10192 21486
rect 10140 21422 10192 21428
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 9772 21072 9824 21078
rect 9678 21040 9734 21049
rect 10152 21049 10180 21422
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 9772 21014 9824 21020
rect 10138 21040 10194 21049
rect 9678 20975 9680 20984
rect 9732 20975 9734 20984
rect 10336 21026 10364 21286
rect 10428 21146 10456 21422
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10138 20975 10194 20984
rect 10232 21004 10284 21010
rect 9680 20946 9732 20952
rect 10336 20998 10456 21026
rect 10520 21010 10548 21927
rect 10612 21554 10640 22510
rect 10876 22432 10928 22438
rect 10876 22374 10928 22380
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10888 21554 10916 22374
rect 11072 21962 11100 22374
rect 11152 22092 11204 22098
rect 11152 22034 11204 22040
rect 11060 21956 11112 21962
rect 11060 21898 11112 21904
rect 10600 21548 10652 21554
rect 10600 21490 10652 21496
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 11072 21486 11100 21898
rect 11164 21486 11192 22034
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 10232 20946 10284 20952
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9600 18902 9628 20742
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9692 19310 9720 20402
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9588 18896 9640 18902
rect 9588 18838 9640 18844
rect 9876 18698 9904 19450
rect 10244 19310 10272 20946
rect 10428 20942 10456 20998
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 10520 19922 10548 20946
rect 10704 20806 10732 21422
rect 11256 21418 11284 21966
rect 11348 21593 11376 22918
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 11980 22704 12032 22710
rect 11980 22646 12032 22652
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11334 21584 11390 21593
rect 11334 21519 11390 21528
rect 11716 21486 11744 22578
rect 11992 22137 12020 22646
rect 11978 22128 12034 22137
rect 11978 22063 12034 22072
rect 12176 22030 12204 22714
rect 12348 22500 12400 22506
rect 12348 22442 12400 22448
rect 12360 22234 12388 22442
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12348 22228 12400 22234
rect 12268 22188 12348 22216
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 12176 21486 12204 21966
rect 12268 21486 12296 22188
rect 12348 22170 12400 22176
rect 12346 22128 12402 22137
rect 12544 22098 12572 22374
rect 12532 22092 12584 22098
rect 12346 22063 12402 22072
rect 12360 21554 12388 22063
rect 12452 22052 12532 22080
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12452 21486 12480 22052
rect 12532 22034 12584 22040
rect 12728 21486 12756 22374
rect 12820 21690 12848 22714
rect 12900 22704 12952 22710
rect 12900 22646 12952 22652
rect 13636 22704 13688 22710
rect 13636 22646 13688 22652
rect 12912 22166 12940 22646
rect 13648 22574 13676 22646
rect 13544 22568 13596 22574
rect 13544 22510 13596 22516
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 13268 22500 13320 22506
rect 13268 22442 13320 22448
rect 13176 22432 13228 22438
rect 13176 22374 13228 22380
rect 12900 22160 12952 22166
rect 12900 22102 12952 22108
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 11704 21480 11756 21486
rect 11704 21422 11756 21428
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 13188 21350 13216 22374
rect 13280 21554 13308 22442
rect 13556 22030 13584 22510
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 13924 22234 13952 22374
rect 13912 22228 13964 22234
rect 13912 22170 13964 22176
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13728 21412 13780 21418
rect 13728 21354 13780 21360
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 11428 21344 11480 21350
rect 11428 21286 11480 21292
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 13176 21344 13228 21350
rect 13176 21286 13228 21292
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13452 21344 13504 21350
rect 13452 21286 13504 21292
rect 13636 21344 13688 21350
rect 13636 21286 13688 21292
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10980 19990 11008 20334
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10508 19916 10560 19922
rect 10508 19858 10560 19864
rect 10980 19310 11008 19926
rect 11164 19922 11192 21286
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10336 18766 10364 19110
rect 10416 18828 10468 18834
rect 10416 18770 10468 18776
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8772 17882 8800 18022
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8864 17626 8892 18022
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 8772 17598 8892 17626
rect 9220 17604 9272 17610
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8680 15502 8708 16934
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 8128 13462 8156 13874
rect 8404 13870 8432 14214
rect 8772 13870 8800 17598
rect 9220 17546 9272 17552
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8864 17134 8892 17478
rect 9232 17134 9260 17546
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 8864 16658 8892 17070
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 9048 16794 9076 17002
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 9232 16658 9260 17070
rect 9416 16726 9444 17818
rect 9784 17814 9812 18566
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9508 17338 9536 17682
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9508 16794 9536 17274
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9784 16538 9812 17750
rect 9876 17678 9904 18634
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9692 16510 9812 16538
rect 9692 16454 9720 16510
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9692 15026 9720 15370
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14550 9720 14758
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8956 13938 8984 14282
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8404 13530 8432 13806
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6840 12714 6868 13262
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6840 12170 6868 12650
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 12374 7420 12582
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5908 11280 5960 11286
rect 5644 11206 5764 11234
rect 5908 11222 5960 11228
rect 5736 11150 5764 11206
rect 6012 11150 6040 11698
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5276 9382 5304 10066
rect 5368 9518 5396 10066
rect 5460 9722 5488 10134
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5552 9518 5580 10066
rect 5644 10062 5672 11018
rect 5736 11014 5764 11086
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5736 10810 5764 10950
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 6012 10724 6040 11086
rect 5920 10696 6040 10724
rect 5920 10606 5948 10696
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 5092 8362 5120 9046
rect 5460 9042 5488 9318
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3252 6934 3280 7278
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3252 6798 3280 6870
rect 3344 6866 3372 7346
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3252 6254 3280 6734
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3344 6186 3372 6802
rect 3436 6458 3464 7142
rect 3620 6730 3648 7482
rect 4080 7478 4108 7686
rect 4172 7546 4200 7686
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 3804 6798 3832 6870
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3608 6724 3660 6730
rect 3608 6666 3660 6672
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3528 5846 3556 6598
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 4080 6458 4108 7278
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4172 6866 4200 7142
rect 4264 7002 4292 7958
rect 4908 7750 4936 8230
rect 5460 7886 5488 8978
rect 5552 8974 5580 9454
rect 6012 9450 6040 9862
rect 6104 9586 6132 10474
rect 6288 10470 6316 11222
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6380 10266 6408 10542
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6380 9654 6408 9930
rect 6564 9722 6592 10066
rect 7024 9926 7052 11018
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5644 8566 5672 8774
rect 6104 8634 6132 8978
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 5632 8560 5684 8566
rect 5684 8520 5764 8548
rect 5632 8502 5684 8508
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4724 6882 4752 7210
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4264 6854 4752 6882
rect 4264 6798 4292 6854
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4172 6254 4200 6666
rect 5092 6254 5120 7686
rect 5460 6798 5488 7822
rect 5644 7546 5672 7958
rect 5736 7954 5764 8520
rect 6380 8498 6408 9590
rect 7116 9110 7144 10474
rect 7208 9518 7236 10678
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7300 10266 7328 10406
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7944 10130 7972 12310
rect 8220 12306 8248 13126
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8404 12374 8432 12718
rect 8496 12434 8524 13398
rect 8588 13394 8616 13806
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8772 13462 8800 13670
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8956 13394 8984 13874
rect 9048 13870 9076 14010
rect 9232 14006 9260 14418
rect 9588 14408 9640 14414
rect 9784 14362 9812 16390
rect 9876 14498 9904 17478
rect 9968 17134 9996 18634
rect 10336 18290 10364 18702
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10428 18222 10456 18770
rect 10888 18766 10916 19246
rect 10980 18902 11008 19246
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 10416 18216 10468 18222
rect 10416 18158 10468 18164
rect 10060 17882 10088 18158
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10244 16998 10272 17070
rect 10888 16998 10916 17070
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10244 16522 10272 16934
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 11440 16046 11468 21286
rect 11612 20528 11664 20534
rect 11612 20470 11664 20476
rect 11624 19310 11652 20470
rect 11992 20398 12020 21286
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12636 20398 12664 20742
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 11992 19378 12020 20334
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12348 19984 12400 19990
rect 12348 19926 12400 19932
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 12084 19310 12112 19858
rect 12164 19440 12216 19446
rect 12164 19382 12216 19388
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 11704 19236 11756 19242
rect 11704 19178 11756 19184
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 9968 14618 9996 15302
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9876 14482 9996 14498
rect 10060 14482 10088 15302
rect 10152 14958 10180 15574
rect 11440 15570 11468 15846
rect 11532 15638 11560 18770
rect 11716 18290 11744 19178
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11796 18692 11848 18698
rect 11796 18634 11848 18640
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11808 17218 11836 18634
rect 11992 18290 12020 18702
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 12084 18222 12112 19246
rect 12176 18834 12204 19382
rect 12268 19310 12296 19858
rect 12360 19378 12388 19926
rect 12544 19378 12572 20198
rect 12636 19922 12664 20334
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 13004 19446 13032 20198
rect 13096 19854 13124 20334
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13096 19514 13124 19790
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12820 18970 12848 19246
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 13004 18766 13032 19382
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 13096 18834 13124 19314
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12900 18148 12952 18154
rect 12900 18090 12952 18096
rect 11716 17190 11836 17218
rect 12912 17202 12940 18090
rect 12900 17196 12952 17202
rect 11716 17134 11744 17190
rect 12900 17138 12952 17144
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11520 15632 11572 15638
rect 11520 15574 11572 15580
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 11244 14952 11296 14958
rect 11440 14906 11468 15506
rect 11624 15502 11652 16050
rect 11716 15910 11744 17070
rect 12912 17066 12940 17138
rect 12900 17060 12952 17066
rect 12900 17002 12952 17008
rect 13372 16658 13400 21286
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13372 16114 13400 16594
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13464 16046 13492 21286
rect 13648 21146 13676 21286
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13740 21010 13768 21354
rect 13832 21010 13860 21966
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13636 20936 13688 20942
rect 13636 20878 13688 20884
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 13556 19310 13584 19722
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13648 17626 13676 20878
rect 13924 19922 13952 21830
rect 14200 21486 14228 21830
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14292 20942 14320 21966
rect 14384 21554 14412 22374
rect 14936 22098 14964 22918
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15108 22228 15160 22234
rect 15108 22170 15160 22176
rect 14924 22092 14976 22098
rect 14924 22034 14976 22040
rect 15120 21690 15148 22170
rect 15212 22030 15240 22714
rect 15304 22506 15332 23054
rect 18144 23044 18196 23050
rect 18144 22986 18196 22992
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 15568 22704 15620 22710
rect 15568 22646 15620 22652
rect 16488 22704 16540 22710
rect 16488 22646 16540 22652
rect 15292 22500 15344 22506
rect 15292 22442 15344 22448
rect 15304 22273 15332 22442
rect 15290 22264 15346 22273
rect 15580 22234 15608 22646
rect 16500 22438 16528 22646
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 15936 22432 15988 22438
rect 15936 22374 15988 22380
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 15290 22199 15346 22208
rect 15568 22228 15620 22234
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 14280 20936 14332 20942
rect 14936 20913 14964 21422
rect 15028 21078 15056 21490
rect 15120 21486 15148 21626
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 15016 21072 15068 21078
rect 15016 21014 15068 21020
rect 15212 21010 15240 21966
rect 15304 21146 15332 22199
rect 15568 22170 15620 22176
rect 15580 21418 15608 22170
rect 15752 22092 15804 22098
rect 15752 22034 15804 22040
rect 15660 22024 15712 22030
rect 15764 22001 15792 22034
rect 15660 21966 15712 21972
rect 15750 21992 15806 22001
rect 15672 21554 15700 21966
rect 15750 21927 15806 21936
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15568 21412 15620 21418
rect 15568 21354 15620 21360
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15396 20942 15424 21354
rect 15948 21010 15976 22374
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 16132 22098 16160 22170
rect 16488 22160 16540 22166
rect 16488 22102 16540 22108
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16212 22092 16264 22098
rect 16212 22034 16264 22040
rect 15936 21004 15988 21010
rect 15936 20946 15988 20952
rect 15384 20936 15436 20942
rect 14280 20878 14332 20884
rect 14922 20904 14978 20913
rect 15384 20878 15436 20884
rect 14922 20839 14978 20848
rect 15948 20058 15976 20946
rect 16224 20874 16252 22034
rect 16500 22001 16528 22102
rect 16486 21992 16542 22001
rect 16486 21927 16542 21936
rect 16592 21010 16620 22510
rect 16684 22506 16712 22918
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17236 22642 17264 22714
rect 17972 22642 18000 22918
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 16672 22500 16724 22506
rect 16672 22442 16724 22448
rect 17132 22500 17184 22506
rect 17132 22442 17184 22448
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 17052 21865 17080 22034
rect 17038 21856 17094 21865
rect 17038 21791 17094 21800
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16684 21146 16712 21422
rect 17052 21418 17080 21791
rect 17144 21622 17172 22442
rect 17132 21616 17184 21622
rect 17132 21558 17184 21564
rect 17040 21412 17092 21418
rect 17040 21354 17092 21360
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 14556 19984 14608 19990
rect 14556 19926 14608 19932
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13832 19242 13860 19654
rect 13924 19378 13952 19858
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13832 18834 13860 19178
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 14016 18766 14044 19314
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14200 19174 14228 19246
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14568 18834 14596 19926
rect 16776 19922 16804 21286
rect 17144 21010 17172 21558
rect 17236 21486 17264 22578
rect 18156 22574 18184 22986
rect 18892 22642 18920 23190
rect 19064 23180 19116 23186
rect 19064 23122 19116 23128
rect 19248 23180 19300 23186
rect 19352 23168 19380 23600
rect 20076 23248 20128 23254
rect 20076 23190 20128 23196
rect 20260 23248 20312 23254
rect 20260 23190 20312 23196
rect 20904 23248 20956 23254
rect 20904 23190 20956 23196
rect 19432 23180 19484 23186
rect 19352 23140 19432 23168
rect 19248 23122 19300 23128
rect 19432 23122 19484 23128
rect 19076 22982 19104 23122
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 19156 22976 19208 22982
rect 19156 22918 19208 22924
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 17316 22500 17368 22506
rect 17316 22442 17368 22448
rect 17328 21690 17356 22442
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 17868 22432 17920 22438
rect 17868 22374 17920 22380
rect 17592 22160 17644 22166
rect 17512 22108 17592 22114
rect 17512 22102 17644 22108
rect 17512 22086 17632 22102
rect 17512 22030 17540 22086
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17696 21894 17724 22374
rect 17774 22264 17830 22273
rect 17774 22199 17830 22208
rect 17788 22098 17816 22199
rect 17776 22092 17828 22098
rect 17776 22034 17828 22040
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17420 21690 17448 21830
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17328 21486 17356 21626
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17224 21480 17276 21486
rect 17224 21422 17276 21428
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17132 21004 17184 21010
rect 17132 20946 17184 20952
rect 17328 20942 17356 21422
rect 17512 21010 17540 21558
rect 17696 21486 17724 21830
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 17316 20936 17368 20942
rect 17316 20878 17368 20884
rect 17788 19990 17816 21490
rect 17880 21146 17908 22374
rect 18800 21894 18828 22510
rect 19076 22098 19104 22918
rect 19168 22642 19196 22918
rect 19260 22710 19288 23122
rect 19248 22704 19300 22710
rect 19248 22646 19300 22652
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 19154 22264 19210 22273
rect 19154 22199 19156 22208
rect 19208 22199 19210 22208
rect 19156 22170 19208 22176
rect 19260 22098 19288 22646
rect 19800 22568 19852 22574
rect 19800 22510 19852 22516
rect 19340 22160 19392 22166
rect 19340 22102 19392 22108
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19352 22030 19380 22102
rect 19340 22024 19392 22030
rect 19812 21978 19840 22510
rect 20088 22438 20116 23190
rect 20168 22976 20220 22982
rect 20168 22918 20220 22924
rect 20180 22574 20208 22918
rect 20272 22574 20300 23190
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20732 22574 20760 22986
rect 20824 22642 20852 23054
rect 20916 22710 20944 23190
rect 22296 23186 22324 23600
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 21192 22982 21220 23122
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 20904 22704 20956 22710
rect 20904 22646 20956 22652
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20168 22568 20220 22574
rect 20168 22510 20220 22516
rect 20260 22568 20312 22574
rect 20260 22510 20312 22516
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 20088 22094 20116 22374
rect 20272 22234 20300 22510
rect 20352 22500 20404 22506
rect 20352 22442 20404 22448
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20364 22166 20392 22442
rect 20824 22166 20852 22578
rect 21192 22574 21220 22918
rect 21468 22778 21496 23122
rect 22652 23112 22704 23118
rect 22652 23054 22704 23060
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21548 22772 21600 22778
rect 21548 22714 21600 22720
rect 21364 22636 21416 22642
rect 21364 22578 21416 22584
rect 21180 22568 21232 22574
rect 21180 22510 21232 22516
rect 21272 22568 21324 22574
rect 21272 22510 21324 22516
rect 21192 22234 21220 22510
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 20352 22160 20404 22166
rect 20350 22128 20352 22137
rect 20812 22160 20864 22166
rect 20404 22128 20406 22137
rect 20168 22094 20220 22098
rect 20088 22092 20220 22094
rect 20088 22066 20168 22092
rect 20812 22102 20864 22108
rect 20350 22063 20406 22072
rect 20168 22034 20220 22040
rect 19340 21966 19392 21972
rect 19720 21962 19840 21978
rect 19708 21956 19840 21962
rect 19760 21950 19840 21956
rect 19708 21898 19760 21904
rect 18696 21888 18748 21894
rect 18788 21888 18840 21894
rect 18696 21830 18748 21836
rect 18786 21856 18788 21865
rect 20536 21888 20588 21894
rect 18840 21856 18842 21865
rect 18708 21690 18736 21830
rect 20536 21830 20588 21836
rect 18786 21791 18842 21800
rect 18696 21684 18748 21690
rect 18696 21626 18748 21632
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 18064 21146 18092 21490
rect 18236 21412 18288 21418
rect 18236 21354 18288 21360
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 18248 21010 18276 21354
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18708 20806 18736 21626
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 20088 21010 20116 21286
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 20364 20874 20392 20946
rect 20352 20868 20404 20874
rect 20352 20810 20404 20816
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19536 20398 19564 20742
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 18972 20324 19024 20330
rect 18972 20266 19024 20272
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 14660 18970 14688 19246
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18290 13952 18566
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 14016 18222 14044 18702
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14200 18426 14228 18566
rect 14292 18426 14320 18770
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 13912 17808 13964 17814
rect 13912 17750 13964 17756
rect 13556 17598 13676 17626
rect 13556 16794 13584 17598
rect 13924 17338 13952 17750
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14568 16794 14596 18226
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 13556 16658 13584 16730
rect 14188 16720 14240 16726
rect 14188 16662 14240 16668
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13556 16182 13584 16594
rect 13740 16250 13768 16594
rect 13728 16244 13780 16250
rect 13648 16204 13728 16232
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 13004 15570 13032 15914
rect 13464 15570 13492 15982
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11520 14952 11572 14958
rect 11296 14900 11520 14906
rect 11244 14894 11572 14900
rect 11256 14878 11560 14894
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10336 14550 10364 14758
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 10600 14544 10652 14550
rect 10652 14504 10732 14532
rect 10600 14486 10652 14492
rect 9864 14476 9996 14482
rect 9916 14470 9996 14476
rect 9864 14418 9916 14424
rect 9588 14350 9640 14356
rect 9600 14074 9628 14350
rect 9692 14334 9812 14362
rect 9968 14362 9996 14470
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9864 14340 9916 14346
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8944 13388 8996 13394
rect 8944 13330 8996 13336
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8496 12406 8616 12434
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8588 12306 8616 12406
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8496 11914 8524 12242
rect 9048 12238 9076 12786
rect 9140 12782 9168 13126
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9232 12306 9260 13942
rect 9692 13818 9720 14334
rect 9968 14334 10088 14362
rect 9864 14282 9916 14288
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9784 13938 9812 14214
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9876 13870 9904 14282
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9864 13864 9916 13870
rect 9600 13802 9720 13818
rect 9588 13796 9720 13802
rect 9640 13790 9720 13796
rect 9862 13832 9864 13841
rect 9916 13832 9918 13841
rect 9862 13767 9918 13776
rect 9588 13738 9640 13744
rect 9968 13394 9996 14214
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 10060 13326 10088 14334
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10152 13870 10180 14214
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10140 13728 10192 13734
rect 10244 13716 10272 14486
rect 10704 14414 10732 14504
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10416 14272 10468 14278
rect 10414 14240 10416 14249
rect 11440 14249 11468 14554
rect 10468 14240 10470 14249
rect 10414 14175 10470 14184
rect 11426 14240 11482 14249
rect 11426 14175 11482 14184
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10324 13864 10376 13870
rect 10428 13852 10456 14010
rect 11440 13870 11468 14175
rect 10376 13824 10456 13852
rect 11060 13864 11112 13870
rect 11058 13832 11060 13841
rect 11428 13864 11480 13870
rect 11112 13832 11114 13841
rect 10324 13806 10376 13812
rect 11428 13806 11480 13812
rect 11058 13767 11114 13776
rect 10192 13688 10272 13716
rect 10140 13670 10192 13676
rect 10244 13394 10272 13688
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 10428 13530 10456 13670
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9324 12782 9352 13126
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9692 12238 9720 12650
rect 9784 12306 9812 13126
rect 11072 12986 11100 13670
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11164 12850 11192 13670
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8496 11898 8616 11914
rect 8496 11892 8628 11898
rect 8496 11886 8576 11892
rect 8576 11834 8628 11840
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8404 11354 8432 11630
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7668 9994 7696 10066
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7484 9518 7512 9862
rect 7852 9722 7880 9862
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 9110 7696 9318
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7546 6592 7686
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6840 7342 6868 8774
rect 7944 8430 7972 8978
rect 8128 8430 8156 9998
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8220 8838 8248 9590
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8312 8974 8340 9522
rect 8496 9382 8524 10134
rect 8588 10062 8616 11834
rect 8680 11694 8708 12038
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8680 10810 8708 11154
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8956 10674 8984 12038
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 10674 9536 10950
rect 9600 10810 9628 11834
rect 10704 11694 10732 12174
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 11286 10732 11630
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 10796 10674 10824 12582
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 10888 10674 10916 12106
rect 10980 11694 11008 12582
rect 11440 12442 11468 12718
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11532 12306 11560 12650
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11716 11898 11744 12174
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 10266 8892 10406
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8864 10062 8892 10202
rect 8956 10130 8984 10474
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8576 10056 8628 10062
rect 8852 10056 8904 10062
rect 8628 10004 8708 10010
rect 8576 9998 8708 10004
rect 8852 9998 8904 10004
rect 8588 9982 8708 9998
rect 8680 9926 8708 9982
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8588 9518 8616 9862
rect 8864 9722 8892 9998
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8956 9586 8984 10066
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7208 8090 7236 8298
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7196 8084 7248 8090
rect 7248 8044 7328 8072
rect 7196 8026 7248 8032
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 6934 5580 7142
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5552 6662 5580 6870
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5736 6322 5764 7210
rect 5828 6866 5856 7210
rect 6012 6866 6040 7210
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 7002 6592 7142
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 5736 5778 5764 6258
rect 5828 6118 5856 6802
rect 6012 6458 6040 6802
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6840 6322 6868 7278
rect 7208 6934 7236 7822
rect 7300 6934 7328 8044
rect 7576 8022 7604 8230
rect 7564 8016 7616 8022
rect 7564 7958 7616 7964
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7576 7002 7604 7754
rect 7852 7750 7880 8230
rect 7944 8022 7972 8366
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7944 7818 7972 7958
rect 8128 7954 8156 8366
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8404 8090 8432 8298
rect 8496 8090 8524 8366
rect 8588 8362 8616 9318
rect 9140 9042 9168 9862
rect 9324 9586 9352 9862
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9416 9382 9444 10134
rect 9508 9518 9536 10610
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 8036 7206 8064 7890
rect 8128 7546 8156 7890
rect 8588 7886 8616 8298
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 8404 6866 8432 7686
rect 8588 7546 8616 7822
rect 8864 7750 8892 8230
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8772 7274 8800 7686
rect 8956 7342 8984 8230
rect 9784 7818 9812 8230
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9876 7410 9904 8434
rect 9956 8016 10008 8022
rect 9954 7984 9956 7993
rect 10324 8016 10376 8022
rect 10008 7984 10010 7993
rect 10324 7958 10376 7964
rect 9954 7919 10010 7928
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8956 6866 8984 7278
rect 9968 6934 9996 7919
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7546 10272 7686
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10244 7002 10272 7210
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 10336 6458 10364 7958
rect 10520 7954 10548 8570
rect 10980 8566 11008 11154
rect 11256 10810 11284 11154
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11440 10130 11468 10746
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11532 10198 11560 10542
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11072 8974 11100 9318
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10888 8430 10916 8502
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10612 7954 10640 8230
rect 10704 8090 10732 8298
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10428 6662 10456 7686
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 10704 6254 10732 8026
rect 10888 6866 10916 8366
rect 10980 7274 11008 8502
rect 11164 8362 11192 8978
rect 11348 8634 11376 9454
rect 11716 8974 11744 9862
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11072 7954 11100 8230
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11164 7936 11192 8298
rect 11348 8090 11376 8570
rect 11808 8430 11836 8978
rect 11900 8430 11928 15098
rect 12084 14958 12112 15370
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12164 14816 12216 14822
rect 12084 14764 12164 14770
rect 12084 14758 12216 14764
rect 12084 14742 12204 14758
rect 12084 14482 12112 14742
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12084 13870 12112 14418
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12440 14068 12492 14074
rect 12360 14028 12440 14056
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12360 13394 12388 14028
rect 12440 14010 12492 14016
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12360 12986 12388 13330
rect 12452 12986 12480 13874
rect 12544 13462 12572 13942
rect 12728 13938 12756 14214
rect 12820 13938 12848 15030
rect 13556 14958 13584 15846
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13188 14482 13216 14758
rect 13556 14482 13584 14894
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12808 13932 12860 13938
rect 12860 13892 12940 13920
rect 12808 13874 12860 13880
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12544 12782 12572 13398
rect 12636 13394 12664 13738
rect 12728 13530 12756 13874
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12820 13530 12848 13670
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 11992 12442 12020 12718
rect 12912 12714 12940 13892
rect 13188 13870 13216 14418
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13280 13394 13308 14350
rect 13556 13870 13584 14418
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13648 13802 13676 16204
rect 13728 16186 13780 16192
rect 14200 16046 14228 16662
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14292 15910 14320 16594
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13728 14952 13780 14958
rect 13832 14940 13860 15438
rect 14292 15162 14320 15846
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 13780 14912 13860 14940
rect 13728 14894 13780 14900
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13740 14482 13768 14758
rect 13728 14476 13780 14482
rect 13832 14464 13860 14912
rect 14476 14618 14504 16594
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 13912 14476 13964 14482
rect 13832 14436 13912 14464
rect 13728 14418 13780 14424
rect 13912 14418 13964 14424
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13740 13530 13768 14418
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 14074 13860 14214
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13832 13938 13860 14010
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13832 13394 13860 13874
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13648 12782 13676 13126
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11992 10606 12020 12378
rect 12268 12374 12296 12582
rect 13556 12434 13584 12718
rect 14016 12442 14044 13262
rect 13464 12406 13584 12434
rect 14004 12436 14056 12442
rect 12256 12368 12308 12374
rect 12256 12310 12308 12316
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12084 10810 12112 11834
rect 13464 11626 13492 12406
rect 14004 12378 14056 12384
rect 14108 11694 14136 13942
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14384 13394 14412 13874
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14384 12434 14412 13330
rect 14660 12442 14688 18226
rect 14752 18222 14780 19450
rect 16868 19378 16896 19722
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 17880 19310 17908 19654
rect 17972 19310 18000 19994
rect 18144 19984 18196 19990
rect 18144 19926 18196 19932
rect 18156 19310 18184 19926
rect 18248 19854 18276 19994
rect 18512 19984 18564 19990
rect 18512 19926 18564 19932
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18248 19310 18276 19654
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 14936 18222 14964 19246
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14936 17202 14964 17682
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 15028 16658 15056 19110
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 15120 18290 15148 18770
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15212 16810 15240 19246
rect 16776 18902 16804 19246
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17144 18902 17172 19110
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 16764 18896 16816 18902
rect 16764 18838 16816 18844
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 16396 18828 16448 18834
rect 16396 18770 16448 18776
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15120 16782 15240 16810
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 15028 16046 15056 16594
rect 15120 16590 15148 16782
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15120 16250 15148 16526
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15120 16114 15148 16186
rect 15212 16182 15240 16594
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15212 15706 15240 15982
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15212 12986 15240 15642
rect 15304 13870 15332 18566
rect 15488 17134 15516 18566
rect 16408 18426 16436 18770
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16500 17746 16528 18566
rect 17604 18222 17632 18566
rect 17696 18222 17724 18906
rect 17972 18290 18000 19110
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17592 18216 17644 18222
rect 17592 18158 17644 18164
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17972 17746 18000 18226
rect 18156 17746 18184 18294
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 18248 17746 18276 18158
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 18144 17740 18196 17746
rect 18144 17682 18196 17688
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 15660 17264 15712 17270
rect 15660 17206 15712 17212
rect 15672 17134 15700 17206
rect 16316 17134 16344 17478
rect 16500 17338 16528 17682
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15396 16658 15424 16934
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15580 16522 15608 16934
rect 15672 16794 15700 17070
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15672 16590 15700 16730
rect 16040 16726 16068 16934
rect 16684 16810 16712 17682
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16776 17134 16804 17478
rect 16868 17134 16896 17614
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17144 17338 17172 17546
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16684 16782 16804 16810
rect 17144 16794 17172 17274
rect 17236 17134 17264 17682
rect 17604 17202 17632 17682
rect 18248 17338 18276 17682
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18340 17338 18368 17478
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18432 17202 18460 18362
rect 18524 17882 18552 19926
rect 18984 19922 19012 20266
rect 19076 19990 19104 20334
rect 19064 19984 19116 19990
rect 19064 19926 19116 19932
rect 19536 19922 19564 20334
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19720 19922 19748 20198
rect 20364 19990 20392 20810
rect 20352 19984 20404 19990
rect 20352 19926 20404 19932
rect 20548 19922 20576 21830
rect 20628 20800 20680 20806
rect 20628 20742 20680 20748
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20640 20602 20668 20742
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20732 20466 20760 20742
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20824 20398 20852 22102
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 21008 21486 21036 21830
rect 21284 21486 21312 22510
rect 21376 22166 21404 22578
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21364 22160 21416 22166
rect 21364 22102 21416 22108
rect 21468 22098 21496 22510
rect 21456 22092 21508 22098
rect 21456 22034 21508 22040
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21008 21078 21036 21286
rect 21284 21146 21312 21286
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 20996 21072 21048 21078
rect 20996 21014 21048 21020
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 21284 20466 21312 20742
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 19524 19916 19576 19922
rect 19524 19858 19576 19864
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 18708 19514 18736 19722
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18880 19304 18932 19310
rect 18880 19246 18932 19252
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 18892 18970 18920 19246
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18788 18216 18840 18222
rect 18892 18204 18920 18906
rect 18972 18216 19024 18222
rect 18892 18176 18972 18204
rect 18788 18158 18840 18164
rect 18972 18158 19024 18164
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18616 17882 18644 18022
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 16672 16720 16724 16726
rect 16672 16662 16724 16668
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 15568 16516 15620 16522
rect 15568 16458 15620 16464
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15396 15910 15424 16390
rect 15672 16114 15700 16526
rect 16212 16516 16264 16522
rect 16212 16458 16264 16464
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 16120 16040 16172 16046
rect 16224 16028 16252 16458
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16316 16250 16344 16390
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16172 16000 16252 16028
rect 16120 15982 16172 15988
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 16224 15570 16252 16000
rect 16316 15910 16344 16050
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15948 14958 15976 15302
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15948 14414 15976 14758
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15488 13530 15516 13738
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15948 13326 15976 14350
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 13462 16068 13670
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14648 12436 14700 12442
rect 14384 12406 14596 12434
rect 14568 12238 14596 12406
rect 14648 12378 14700 12384
rect 14936 12306 14964 12582
rect 16224 12374 16252 15506
rect 16408 14890 16436 16526
rect 16684 16182 16712 16662
rect 16776 16250 16804 16782
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 18064 16522 18092 17070
rect 18524 16794 18552 17070
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18052 16516 18104 16522
rect 18052 16458 18104 16464
rect 18616 16250 18644 17818
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18708 17134 18736 17682
rect 18800 17542 18828 18158
rect 19168 17746 19196 19246
rect 19536 19242 19564 19654
rect 19524 19236 19576 19242
rect 19524 19178 19576 19184
rect 19996 18970 20024 19790
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19720 18222 19748 18770
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18708 16658 18736 17070
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16776 16046 16804 16186
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16500 15638 16528 15982
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16592 15638 16620 15846
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16684 15570 16712 15846
rect 16960 15570 16988 16118
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 16776 14550 16804 15302
rect 16868 15162 16896 15438
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 16764 14544 16816 14550
rect 16764 14486 16816 14492
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16776 13530 16804 14010
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 16316 12306 16344 13262
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14568 11898 14596 12174
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14660 11694 14688 12038
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 13464 11218 13492 11562
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 11286 13860 11494
rect 14292 11354 14320 11630
rect 14936 11354 14964 12242
rect 15120 11898 15148 12242
rect 16408 12238 16436 13330
rect 17052 13326 17080 15098
rect 17144 13938 17172 15302
rect 17328 14958 17356 15506
rect 18800 15366 18828 17478
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19260 16658 19288 16934
rect 19720 16726 19748 18158
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 19904 17814 19932 18022
rect 19892 17808 19944 17814
rect 19892 17750 19944 17756
rect 19708 16720 19760 16726
rect 19708 16662 19760 16668
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 16046 19288 16594
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19444 16114 19472 16186
rect 19524 16176 19576 16182
rect 19708 16176 19760 16182
rect 19576 16124 19708 16130
rect 19524 16118 19760 16124
rect 19432 16108 19484 16114
rect 19536 16102 19748 16118
rect 19432 16050 19484 16056
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 17328 14618 17356 14894
rect 17776 14884 17828 14890
rect 17776 14826 17828 14832
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17788 14482 17816 14826
rect 17972 14618 18000 14894
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17788 14006 17816 14418
rect 18064 14278 18092 14894
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18340 14550 18368 14826
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17788 13870 17816 13942
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17144 13530 17172 13670
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 14280 11348 14332 11354
rect 14924 11348 14976 11354
rect 14280 11290 14332 11296
rect 14844 11308 14924 11336
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 12360 10606 12388 10950
rect 14292 10810 14320 11290
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 12084 10130 12112 10474
rect 12360 10266 12388 10542
rect 12452 10470 12480 10678
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12820 10130 12848 10406
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12360 9586 12388 9862
rect 13648 9586 13676 10406
rect 14200 10062 14228 10406
rect 14292 10130 14320 10746
rect 14844 10606 14872 11308
rect 14924 11290 14976 11296
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14936 10674 14964 11154
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 10130 14780 10406
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14924 9988 14976 9994
rect 14924 9930 14976 9936
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14476 9586 14504 9862
rect 14936 9586 14964 9930
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12268 8838 12296 9318
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11532 8090 11560 8366
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11244 7948 11296 7954
rect 11164 7908 11244 7936
rect 11164 7818 11192 7908
rect 11244 7890 11296 7896
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11244 7540 11296 7546
rect 11348 7528 11376 8026
rect 11532 7546 11560 8026
rect 11624 7954 11652 8230
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11296 7500 11376 7528
rect 11520 7540 11572 7546
rect 11244 7482 11296 7488
rect 11520 7482 11572 7488
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10980 6866 11008 7210
rect 11072 6866 11100 7482
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 11624 6186 11652 7890
rect 11716 7206 11744 7958
rect 11808 7750 11836 8230
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11900 7206 11928 8366
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 12360 7002 12388 8298
rect 12716 8016 12768 8022
rect 12714 7984 12716 7993
rect 12768 7984 12770 7993
rect 13004 7954 13032 8434
rect 13740 8362 13768 9454
rect 14384 9042 14412 9454
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14384 8634 14412 8978
rect 15028 8974 15056 11562
rect 15120 11218 15148 11834
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15120 10606 15148 11154
rect 16224 10606 16252 11222
rect 16408 11082 16436 12174
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16408 10606 16436 11018
rect 16592 10656 16620 11154
rect 16684 11150 16712 12038
rect 16960 11218 16988 12242
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16592 10628 16712 10656
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16592 9654 16620 10474
rect 16684 9994 16712 10628
rect 16868 10606 16896 10950
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16684 9722 16712 9930
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16684 9518 16712 9658
rect 15200 9512 15252 9518
rect 16672 9512 16724 9518
rect 15200 9454 15252 9460
rect 16486 9480 16542 9489
rect 15212 9110 15240 9454
rect 15476 9444 15528 9450
rect 16672 9454 16724 9460
rect 16486 9415 16542 9424
rect 16764 9444 16816 9450
rect 15476 9386 15528 9392
rect 15488 9178 15516 9386
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 16500 9110 16528 9415
rect 16764 9386 16816 9392
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 14556 8968 14608 8974
rect 15016 8968 15068 8974
rect 14556 8910 14608 8916
rect 14936 8916 15016 8922
rect 14936 8910 15068 8916
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13096 8090 13124 8298
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 12714 7919 12770 7928
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12452 7342 12480 7686
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 13004 6866 13032 7890
rect 13188 7546 13216 8230
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13372 7342 13400 7686
rect 13464 7478 13492 8230
rect 13924 8090 13952 8570
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14292 8090 14320 8230
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14384 7954 14412 8570
rect 14476 8362 14504 8842
rect 14568 8498 14596 8910
rect 14936 8894 15056 8910
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14568 8362 14596 8434
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14476 7546 14504 8298
rect 14660 8022 14688 8502
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 7002 13216 7142
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13556 6934 13584 7482
rect 14752 7342 14780 8230
rect 14936 7954 14964 8894
rect 15212 8566 15240 9046
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 15028 8090 15056 8298
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 14936 7750 14964 7890
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 15212 7342 15240 8502
rect 16316 8498 16344 8910
rect 16592 8906 16620 9318
rect 16776 9178 16804 9386
rect 16868 9382 16896 10406
rect 16960 10130 16988 11154
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17052 10810 17080 10950
rect 17236 10810 17264 13738
rect 17868 13388 17920 13394
rect 17972 13376 18000 13942
rect 18064 13462 18092 14010
rect 18248 13870 18276 14214
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 18340 13394 18368 14486
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 18420 13456 18472 13462
rect 18420 13398 18472 13404
rect 17920 13348 18000 13376
rect 18328 13388 18380 13394
rect 17868 13330 17920 13336
rect 18328 13330 18380 13336
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18064 12714 18092 13262
rect 18432 12918 18460 13398
rect 18524 13190 18552 14418
rect 18616 14414 18644 14962
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18708 13802 18736 15098
rect 19168 15026 19196 15982
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19260 14958 19288 15982
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 19536 15570 19564 15846
rect 19720 15570 19748 15846
rect 20180 15706 20208 19858
rect 20640 19174 20668 20334
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20732 19718 20760 19858
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20628 19168 20680 19174
rect 20628 19110 20680 19116
rect 20364 18834 20392 19110
rect 20640 18834 20668 19110
rect 20352 18828 20404 18834
rect 20352 18770 20404 18776
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20364 16046 20392 18770
rect 20732 17542 20760 19654
rect 20916 17746 20944 20198
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21100 19310 21128 19654
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21192 19242 21220 19926
rect 21284 19854 21312 20402
rect 21468 20398 21496 22034
rect 21560 21622 21588 22714
rect 21652 22642 21680 22918
rect 21824 22704 21876 22710
rect 21824 22646 21876 22652
rect 21640 22636 21692 22642
rect 21640 22578 21692 22584
rect 21652 21962 21680 22578
rect 21836 22094 21864 22646
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22112 22234 22140 22374
rect 22100 22228 22152 22234
rect 22100 22170 22152 22176
rect 22204 22098 22232 22374
rect 22664 22166 22692 23054
rect 22652 22160 22704 22166
rect 22374 22128 22430 22137
rect 21744 22066 21864 22094
rect 22192 22092 22244 22098
rect 21744 22030 21772 22066
rect 22652 22102 22704 22108
rect 22374 22063 22376 22072
rect 22192 22034 22244 22040
rect 22428 22063 22430 22072
rect 22376 22034 22428 22040
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 21640 21956 21692 21962
rect 21640 21898 21692 21904
rect 21744 21690 21772 21966
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 21548 21616 21600 21622
rect 21548 21558 21600 21564
rect 21560 21078 21588 21558
rect 22296 21554 22324 21966
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 22296 21010 22324 21490
rect 22284 21004 22336 21010
rect 22284 20946 22336 20952
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 22652 20392 22704 20398
rect 22652 20334 22704 20340
rect 21468 20058 21496 20334
rect 21824 20324 21876 20330
rect 21824 20266 21876 20272
rect 22468 20324 22520 20330
rect 22468 20266 22520 20272
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 21100 17338 21128 18770
rect 21192 18766 21220 19178
rect 21836 18970 21864 20266
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 22008 20256 22060 20262
rect 22008 20198 22060 20204
rect 21928 19854 21956 20198
rect 22020 19990 22048 20198
rect 22008 19984 22060 19990
rect 22008 19926 22060 19932
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22204 19514 22232 19654
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 21192 17678 21220 18702
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21376 18222 21404 18566
rect 21916 18420 21968 18426
rect 21916 18362 21968 18368
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 21364 18216 21416 18222
rect 21284 18176 21364 18204
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 20812 15972 20864 15978
rect 20812 15914 20864 15920
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 20732 15570 20760 15846
rect 20824 15706 20852 15914
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19708 15564 19760 15570
rect 19708 15506 19760 15512
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20824 15434 20852 15642
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 19720 15026 19748 15302
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 20548 14958 20576 15302
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 20444 14952 20496 14958
rect 20444 14894 20496 14900
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19444 14618 19472 14826
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18696 13796 18748 13802
rect 18696 13738 18748 13744
rect 18800 13530 18828 14350
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17972 12374 18000 12582
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 17328 11354 17356 12310
rect 17788 11898 17816 12310
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 18064 11694 18092 12310
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18432 11626 18460 12854
rect 18524 12782 18552 13126
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18420 11620 18472 11626
rect 18420 11562 18472 11568
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17236 10266 17264 10746
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 17328 9178 17356 11290
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17788 10538 17816 11222
rect 18432 11218 18460 11562
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17420 9518 17448 10066
rect 17604 9994 17632 10202
rect 17788 10130 17816 10474
rect 17880 10266 17908 10950
rect 18248 10606 18276 10950
rect 18708 10674 18736 12174
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17420 9110 17448 9454
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 17408 9104 17460 9110
rect 17408 9046 17460 9052
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16500 8430 16528 8774
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16500 8022 16528 8366
rect 16684 8090 16712 9046
rect 17420 8498 17448 9046
rect 17604 8838 17632 9930
rect 17788 9110 17816 10066
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17788 8634 17816 9046
rect 17880 8906 17908 10066
rect 18708 9586 18736 10610
rect 18984 10470 19012 14418
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 19076 14074 19104 14214
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19076 12442 19104 12718
rect 19168 12646 19196 13330
rect 20456 13326 20484 14894
rect 20732 13410 20760 15302
rect 20916 15026 20944 17274
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 21008 15162 21036 15302
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 21284 14074 21312 18176
rect 21364 18158 21416 18164
rect 21732 18216 21784 18222
rect 21732 18158 21784 18164
rect 21744 18034 21772 18158
rect 21928 18154 21956 18362
rect 21916 18148 21968 18154
rect 21916 18090 21968 18096
rect 22020 18034 22048 18362
rect 21744 18006 22048 18034
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 21548 17536 21600 17542
rect 21548 17478 21600 17484
rect 21560 16658 21588 17478
rect 22020 17338 22048 17682
rect 22008 17332 22060 17338
rect 22008 17274 22060 17280
rect 21824 16720 21876 16726
rect 21824 16662 21876 16668
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21560 16250 21588 16594
rect 21640 16448 21692 16454
rect 21640 16390 21692 16396
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21468 15026 21496 16050
rect 21652 16046 21680 16390
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21652 15502 21680 15846
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20548 13382 20760 13410
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20548 13326 20576 13382
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19352 12714 19380 13194
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 19720 12782 19748 13126
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 12442 19196 12582
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19168 11694 19196 12378
rect 19444 12102 19472 12718
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19444 11830 19472 12038
rect 19812 11898 19840 13126
rect 20456 12986 20484 13262
rect 20640 13190 20668 13262
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19432 11824 19484 11830
rect 19432 11766 19484 11772
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19444 11218 19472 11766
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18064 8974 18092 9522
rect 19156 9444 19208 9450
rect 19156 9386 19208 9392
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18800 9110 18828 9318
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17788 8430 17816 8570
rect 18616 8514 18644 8978
rect 18616 8498 18736 8514
rect 18616 8492 18748 8498
rect 18616 8486 18696 8492
rect 18696 8434 18748 8440
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 19168 8412 19196 9386
rect 19444 9110 19472 11154
rect 19720 10810 19748 11154
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19996 10538 20024 11494
rect 20180 11354 20208 12038
rect 20272 11626 20300 12242
rect 20456 12238 20484 12922
rect 20640 12374 20668 13126
rect 20732 12782 20760 13382
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20456 11694 20484 12174
rect 20732 11694 20760 12718
rect 20824 12646 20852 13398
rect 20916 12986 20944 13806
rect 21376 13734 21404 14894
rect 21652 14414 21680 15438
rect 21836 14618 21864 16662
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 22112 16250 22140 16526
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22204 16114 22232 19450
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22296 18902 22324 19110
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22388 18834 22416 19858
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22480 18630 22508 20266
rect 22664 19310 22692 20334
rect 22744 19916 22796 19922
rect 22744 19858 22796 19864
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22560 19236 22612 19242
rect 22560 19178 22612 19184
rect 22572 18970 22600 19178
rect 22560 18964 22612 18970
rect 22560 18906 22612 18912
rect 22468 18624 22520 18630
rect 22468 18566 22520 18572
rect 22572 16590 22600 18906
rect 22756 18306 22784 19858
rect 22836 19848 22888 19854
rect 22836 19790 22888 19796
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 22848 19310 22876 19790
rect 23032 19689 23060 19790
rect 23018 19680 23074 19689
rect 23018 19615 23074 19624
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 22940 18426 22968 18770
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 22928 18420 22980 18426
rect 22928 18362 22980 18368
rect 22664 18278 22784 18306
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22664 16250 22692 18278
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22756 17882 22784 18158
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22848 17746 22876 18362
rect 22928 18080 22980 18086
rect 23032 18034 23060 18566
rect 22980 18028 23060 18034
rect 22928 18022 23060 18028
rect 22940 18006 23060 18022
rect 23032 17746 23060 18006
rect 22836 17740 22888 17746
rect 22836 17682 22888 17688
rect 23020 17740 23072 17746
rect 23020 17682 23072 17688
rect 22744 17060 22796 17066
rect 22744 17002 22796 17008
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22204 15570 22232 16050
rect 22192 15564 22244 15570
rect 22192 15506 22244 15512
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 22112 14958 22140 15302
rect 22664 15042 22692 16186
rect 22572 15014 22692 15042
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21836 14482 21864 14554
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21744 14362 21772 14418
rect 22020 14362 22048 14418
rect 21744 14334 22048 14362
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 13394 21404 13670
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 21272 13252 21324 13258
rect 21272 13194 21324 13200
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 21008 12714 21036 13194
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 12986 21128 13126
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 20996 12708 21048 12714
rect 20996 12650 21048 12656
rect 20812 12640 20864 12646
rect 20864 12600 20944 12628
rect 20812 12582 20864 12588
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20720 11688 20772 11694
rect 20772 11636 20852 11642
rect 20720 11630 20852 11636
rect 20260 11620 20312 11626
rect 20732 11614 20852 11630
rect 20260 11562 20312 11568
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20180 10538 20208 11290
rect 20732 10810 20760 11494
rect 20824 11354 20852 11614
rect 20916 11540 20944 12600
rect 21008 12442 21036 12650
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 21008 11762 21036 12378
rect 21284 11898 21312 13194
rect 21376 12986 21404 13330
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21560 12764 21588 14010
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21376 12736 21588 12764
rect 21376 12434 21404 12736
rect 21652 12442 21680 13330
rect 21640 12436 21692 12442
rect 21376 12406 21588 12434
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 20996 11552 21048 11558
rect 20916 11512 20996 11540
rect 20996 11494 21048 11500
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 21008 11150 21036 11494
rect 20996 11144 21048 11150
rect 20996 11086 21048 11092
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 19984 10532 20036 10538
rect 19984 10474 20036 10480
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 20824 10248 20852 11018
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20640 10220 20852 10248
rect 20640 9602 20668 10220
rect 20916 10130 20944 10746
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20732 9722 20760 10066
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20640 9574 20760 9602
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19248 8424 19300 8430
rect 19168 8384 19248 8412
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16500 7818 16528 7958
rect 16960 7818 16988 8298
rect 17788 7954 17816 8366
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 17972 7750 18000 8230
rect 18156 8022 18184 8230
rect 18800 8090 18828 8298
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18144 8016 18196 8022
rect 18144 7958 18196 7964
rect 19168 7750 19196 8384
rect 19248 8366 19300 8372
rect 19432 8356 19484 8362
rect 19432 8298 19484 8304
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 15396 7546 15424 7686
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 19444 7342 19472 8298
rect 19536 8090 19564 9318
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19628 7970 19656 9386
rect 19904 9178 19932 9386
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19536 7954 19656 7970
rect 19524 7948 19656 7954
rect 19576 7942 19656 7948
rect 19524 7890 19576 7896
rect 19536 7546 19564 7890
rect 19720 7886 19748 8978
rect 19904 8090 19932 9114
rect 20076 8968 20128 8974
rect 20364 8945 20392 9114
rect 20076 8910 20128 8916
rect 20350 8936 20406 8945
rect 20088 8634 20116 8910
rect 20350 8871 20406 8880
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 20088 7410 20116 8570
rect 20168 8288 20220 8294
rect 20168 8230 20220 8236
rect 20180 8022 20208 8230
rect 20168 8016 20220 8022
rect 20168 7958 20220 7964
rect 20732 7750 20760 9574
rect 20824 9450 20852 9930
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20916 9178 20944 10066
rect 21008 9364 21036 11086
rect 21100 10538 21128 11630
rect 21376 11082 21404 12310
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21088 10532 21140 10538
rect 21088 10474 21140 10480
rect 21100 10198 21128 10474
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 21100 9518 21128 10134
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 21192 9586 21220 10066
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 21088 9376 21140 9382
rect 21008 9336 21088 9364
rect 21088 9318 21140 9324
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20824 8838 20852 8978
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20824 8498 20852 8774
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20824 8090 20852 8434
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20916 7342 20944 8570
rect 21008 8430 21036 9046
rect 21100 8634 21128 9318
rect 21180 9036 21232 9042
rect 21180 8978 21232 8984
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 21008 8022 21036 8366
rect 21192 8294 21220 8978
rect 21284 8294 21312 9862
rect 21376 9722 21404 9862
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21364 9512 21416 9518
rect 21362 9480 21364 9489
rect 21416 9480 21418 9489
rect 21362 9415 21418 9424
rect 21468 9178 21496 9998
rect 21560 9518 21588 12406
rect 21640 12378 21692 12384
rect 21652 11354 21680 12378
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21744 11218 21772 13466
rect 21836 12850 21864 13670
rect 22020 13394 22048 14334
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 22008 13388 22060 13394
rect 22008 13330 22060 13336
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 21928 11014 21956 13126
rect 22112 12714 22140 13398
rect 22100 12708 22152 12714
rect 22100 12650 22152 12656
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 22020 11354 22048 12242
rect 22112 11354 22140 12650
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 21916 11008 21968 11014
rect 21916 10950 21968 10956
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 21732 10736 21784 10742
rect 21732 10678 21784 10684
rect 21640 10532 21692 10538
rect 21640 10474 21692 10480
rect 21652 10130 21680 10474
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21744 9738 21772 10678
rect 22020 10198 22048 10950
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22112 10266 22140 10406
rect 22204 10266 22232 14418
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22296 14090 22324 14350
rect 22388 14278 22416 14758
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22376 14272 22428 14278
rect 22376 14214 22428 14220
rect 22296 14062 22416 14090
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22296 12374 22324 12718
rect 22284 12368 22336 12374
rect 22284 12310 22336 12316
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22296 11014 22324 11494
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22008 10192 22060 10198
rect 22008 10134 22060 10140
rect 22388 9926 22416 14062
rect 22480 10470 22508 14418
rect 22572 14414 22600 15014
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 22664 13394 22692 14894
rect 22756 13938 22784 17002
rect 22848 14618 22876 17682
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 22848 14006 22876 14554
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22664 11558 22692 13330
rect 22756 12434 22784 13874
rect 22756 12406 22876 12434
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22848 10810 22876 12406
rect 23018 11792 23074 11801
rect 23018 11727 23074 11736
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22572 9926 22600 10746
rect 23032 10606 23060 11727
rect 23020 10600 23072 10606
rect 23020 10542 23072 10548
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22560 9920 22612 9926
rect 22560 9862 22612 9868
rect 21652 9710 21772 9738
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 21456 9172 21508 9178
rect 21456 9114 21508 9120
rect 21652 8430 21680 9710
rect 21824 9444 21876 9450
rect 21824 9386 21876 9392
rect 21640 8424 21692 8430
rect 21640 8366 21692 8372
rect 21652 8294 21680 8366
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 20996 8016 21048 8022
rect 20996 7958 21048 7964
rect 21100 7342 21128 8230
rect 21364 8016 21416 8022
rect 21364 7958 21416 7964
rect 21376 7342 21404 7958
rect 21548 7948 21600 7954
rect 21548 7890 21600 7896
rect 21560 7546 21588 7890
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 21652 7410 21680 8230
rect 21836 7954 21864 9386
rect 22572 9178 22600 9862
rect 22560 9172 22612 9178
rect 22560 9114 22612 9120
rect 22756 8945 22784 10066
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 22848 9722 22876 9998
rect 22836 9716 22888 9722
rect 22836 9658 22888 9664
rect 22742 8936 22798 8945
rect 22742 8871 22798 8880
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 21916 8356 21968 8362
rect 21916 8298 21968 8304
rect 21928 8090 21956 8298
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 22020 8022 22048 8774
rect 22652 8356 22704 8362
rect 22652 8298 22704 8304
rect 22664 8090 22692 8298
rect 22652 8084 22704 8090
rect 22652 8026 22704 8032
rect 22008 8016 22060 8022
rect 22008 7958 22060 7964
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 21836 7546 21864 7890
rect 22020 7750 22048 7958
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 21088 7336 21140 7342
rect 21088 7278 21140 7284
rect 21364 7336 21416 7342
rect 21364 7278 21416 7284
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5828 5914 5856 6054
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 22756 4146 22784 7278
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22928 4004 22980 4010
rect 22928 3946 22980 3952
rect 22940 3913 22968 3946
rect 22926 3904 22982 3913
rect 4322 3836 4630 3845
rect 22926 3839 22982 3848
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
<< via2 >>
rect 4328 23418 4384 23420
rect 4408 23418 4464 23420
rect 4488 23418 4544 23420
rect 4568 23418 4624 23420
rect 4328 23366 4374 23418
rect 4374 23366 4384 23418
rect 4408 23366 4438 23418
rect 4438 23366 4450 23418
rect 4450 23366 4464 23418
rect 4488 23366 4502 23418
rect 4502 23366 4514 23418
rect 4514 23366 4544 23418
rect 4568 23366 4578 23418
rect 4578 23366 4624 23418
rect 4328 23364 4384 23366
rect 4408 23364 4464 23366
rect 4488 23364 4544 23366
rect 4568 23364 4624 23366
rect 3668 22874 3724 22876
rect 3748 22874 3804 22876
rect 3828 22874 3884 22876
rect 3908 22874 3964 22876
rect 3668 22822 3714 22874
rect 3714 22822 3724 22874
rect 3748 22822 3778 22874
rect 3778 22822 3790 22874
rect 3790 22822 3804 22874
rect 3828 22822 3842 22874
rect 3842 22822 3854 22874
rect 3854 22822 3884 22874
rect 3908 22822 3918 22874
rect 3918 22822 3964 22874
rect 3668 22820 3724 22822
rect 3748 22820 3804 22822
rect 3828 22820 3884 22822
rect 3908 22820 3964 22822
rect 4328 22330 4384 22332
rect 4408 22330 4464 22332
rect 4488 22330 4544 22332
rect 4568 22330 4624 22332
rect 4328 22278 4374 22330
rect 4374 22278 4384 22330
rect 4408 22278 4438 22330
rect 4438 22278 4450 22330
rect 4450 22278 4464 22330
rect 4488 22278 4502 22330
rect 4502 22278 4514 22330
rect 4514 22278 4544 22330
rect 4568 22278 4578 22330
rect 4578 22278 4624 22330
rect 4328 22276 4384 22278
rect 4408 22276 4464 22278
rect 4488 22276 4544 22278
rect 4568 22276 4624 22278
rect 3668 21786 3724 21788
rect 3748 21786 3804 21788
rect 3828 21786 3884 21788
rect 3908 21786 3964 21788
rect 3668 21734 3714 21786
rect 3714 21734 3724 21786
rect 3748 21734 3778 21786
rect 3778 21734 3790 21786
rect 3790 21734 3804 21786
rect 3828 21734 3842 21786
rect 3842 21734 3854 21786
rect 3854 21734 3884 21786
rect 3908 21734 3918 21786
rect 3918 21734 3964 21786
rect 3668 21732 3724 21734
rect 3748 21732 3804 21734
rect 3828 21732 3884 21734
rect 3908 21732 3964 21734
rect 3668 20698 3724 20700
rect 3748 20698 3804 20700
rect 3828 20698 3884 20700
rect 3908 20698 3964 20700
rect 3668 20646 3714 20698
rect 3714 20646 3724 20698
rect 3748 20646 3778 20698
rect 3778 20646 3790 20698
rect 3790 20646 3804 20698
rect 3828 20646 3842 20698
rect 3842 20646 3854 20698
rect 3854 20646 3884 20698
rect 3908 20646 3918 20698
rect 3918 20646 3964 20698
rect 3668 20644 3724 20646
rect 3748 20644 3804 20646
rect 3828 20644 3884 20646
rect 3908 20644 3964 20646
rect 4328 21242 4384 21244
rect 4408 21242 4464 21244
rect 4488 21242 4544 21244
rect 4568 21242 4624 21244
rect 4328 21190 4374 21242
rect 4374 21190 4384 21242
rect 4408 21190 4438 21242
rect 4438 21190 4450 21242
rect 4450 21190 4464 21242
rect 4488 21190 4502 21242
rect 4502 21190 4514 21242
rect 4514 21190 4544 21242
rect 4568 21190 4578 21242
rect 4578 21190 4624 21242
rect 4328 21188 4384 21190
rect 4408 21188 4464 21190
rect 4488 21188 4544 21190
rect 4568 21188 4624 21190
rect 3668 19610 3724 19612
rect 3748 19610 3804 19612
rect 3828 19610 3884 19612
rect 3908 19610 3964 19612
rect 3668 19558 3714 19610
rect 3714 19558 3724 19610
rect 3748 19558 3778 19610
rect 3778 19558 3790 19610
rect 3790 19558 3804 19610
rect 3828 19558 3842 19610
rect 3842 19558 3854 19610
rect 3854 19558 3884 19610
rect 3908 19558 3918 19610
rect 3918 19558 3964 19610
rect 3668 19556 3724 19558
rect 3748 19556 3804 19558
rect 3828 19556 3884 19558
rect 3908 19556 3964 19558
rect 4328 20154 4384 20156
rect 4408 20154 4464 20156
rect 4488 20154 4544 20156
rect 4568 20154 4624 20156
rect 4328 20102 4374 20154
rect 4374 20102 4384 20154
rect 4408 20102 4438 20154
rect 4438 20102 4450 20154
rect 4450 20102 4464 20154
rect 4488 20102 4502 20154
rect 4502 20102 4514 20154
rect 4514 20102 4544 20154
rect 4568 20102 4578 20154
rect 4578 20102 4624 20154
rect 4328 20100 4384 20102
rect 4408 20100 4464 20102
rect 4488 20100 4544 20102
rect 4568 20100 4624 20102
rect 4802 19252 4804 19272
rect 4804 19252 4856 19272
rect 4856 19252 4858 19272
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 4802 19216 4858 19252
rect 4328 19066 4384 19068
rect 4408 19066 4464 19068
rect 4488 19066 4544 19068
rect 4568 19066 4624 19068
rect 4328 19014 4374 19066
rect 4374 19014 4384 19066
rect 4408 19014 4438 19066
rect 4438 19014 4450 19066
rect 4450 19014 4464 19066
rect 4488 19014 4502 19066
rect 4502 19014 4514 19066
rect 4514 19014 4544 19066
rect 4568 19014 4578 19066
rect 4578 19014 4624 19066
rect 4328 19012 4384 19014
rect 4408 19012 4464 19014
rect 4488 19012 4544 19014
rect 4568 19012 4624 19014
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 4328 17978 4384 17980
rect 4408 17978 4464 17980
rect 4488 17978 4544 17980
rect 4568 17978 4624 17980
rect 4328 17926 4374 17978
rect 4374 17926 4384 17978
rect 4408 17926 4438 17978
rect 4438 17926 4450 17978
rect 4450 17926 4464 17978
rect 4488 17926 4502 17978
rect 4502 17926 4514 17978
rect 4514 17926 4544 17978
rect 4568 17926 4578 17978
rect 4578 17926 4624 17978
rect 4328 17924 4384 17926
rect 4408 17924 4464 17926
rect 4488 17924 4544 17926
rect 4568 17924 4624 17926
rect 4328 16890 4384 16892
rect 4408 16890 4464 16892
rect 4488 16890 4544 16892
rect 4568 16890 4624 16892
rect 4328 16838 4374 16890
rect 4374 16838 4384 16890
rect 4408 16838 4438 16890
rect 4438 16838 4450 16890
rect 4450 16838 4464 16890
rect 4488 16838 4502 16890
rect 4502 16838 4514 16890
rect 4514 16838 4544 16890
rect 4568 16838 4578 16890
rect 4578 16838 4624 16890
rect 4328 16836 4384 16838
rect 4408 16836 4464 16838
rect 4488 16836 4544 16838
rect 4568 16836 4624 16838
rect 4328 15802 4384 15804
rect 4408 15802 4464 15804
rect 4488 15802 4544 15804
rect 4568 15802 4624 15804
rect 4328 15750 4374 15802
rect 4374 15750 4384 15802
rect 4408 15750 4438 15802
rect 4438 15750 4450 15802
rect 4450 15750 4464 15802
rect 4488 15750 4502 15802
rect 4502 15750 4514 15802
rect 4514 15750 4544 15802
rect 4568 15750 4578 15802
rect 4578 15750 4624 15802
rect 4328 15748 4384 15750
rect 4408 15748 4464 15750
rect 4488 15748 4544 15750
rect 4568 15748 4624 15750
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 6090 20848 6146 20904
rect 5538 19216 5594 19272
rect 4328 14714 4384 14716
rect 4408 14714 4464 14716
rect 4488 14714 4544 14716
rect 4568 14714 4624 14716
rect 4328 14662 4374 14714
rect 4374 14662 4384 14714
rect 4408 14662 4438 14714
rect 4438 14662 4450 14714
rect 4450 14662 4464 14714
rect 4488 14662 4502 14714
rect 4502 14662 4514 14714
rect 4514 14662 4544 14714
rect 4568 14662 4578 14714
rect 4578 14662 4624 14714
rect 4328 14660 4384 14662
rect 4408 14660 4464 14662
rect 4488 14660 4544 14662
rect 4568 14660 4624 14662
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 4328 13626 4384 13628
rect 4408 13626 4464 13628
rect 4488 13626 4544 13628
rect 4568 13626 4624 13628
rect 4328 13574 4374 13626
rect 4374 13574 4384 13626
rect 4408 13574 4438 13626
rect 4438 13574 4450 13626
rect 4450 13574 4464 13626
rect 4488 13574 4502 13626
rect 4502 13574 4514 13626
rect 4514 13574 4544 13626
rect 4568 13574 4578 13626
rect 4578 13574 4624 13626
rect 4328 13572 4384 13574
rect 4408 13572 4464 13574
rect 4488 13572 4544 13574
rect 4568 13572 4624 13574
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 4328 12538 4384 12540
rect 4408 12538 4464 12540
rect 4488 12538 4544 12540
rect 4568 12538 4624 12540
rect 4328 12486 4374 12538
rect 4374 12486 4384 12538
rect 4408 12486 4438 12538
rect 4438 12486 4450 12538
rect 4450 12486 4464 12538
rect 4488 12486 4502 12538
rect 4502 12486 4514 12538
rect 4514 12486 4544 12538
rect 4568 12486 4578 12538
rect 4578 12486 4624 12538
rect 4328 12484 4384 12486
rect 4408 12484 4464 12486
rect 4488 12484 4544 12486
rect 4568 12484 4624 12486
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 5354 13640 5410 13696
rect 4328 11450 4384 11452
rect 4408 11450 4464 11452
rect 4488 11450 4544 11452
rect 4568 11450 4624 11452
rect 4328 11398 4374 11450
rect 4374 11398 4384 11450
rect 4408 11398 4438 11450
rect 4438 11398 4450 11450
rect 4450 11398 4464 11450
rect 4488 11398 4502 11450
rect 4502 11398 4514 11450
rect 4514 11398 4544 11450
rect 4568 11398 4578 11450
rect 4578 11398 4624 11450
rect 4328 11396 4384 11398
rect 4408 11396 4464 11398
rect 4488 11396 4544 11398
rect 4568 11396 4624 11398
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 4328 10362 4384 10364
rect 4408 10362 4464 10364
rect 4488 10362 4544 10364
rect 4568 10362 4624 10364
rect 4328 10310 4374 10362
rect 4374 10310 4384 10362
rect 4408 10310 4438 10362
rect 4438 10310 4450 10362
rect 4450 10310 4464 10362
rect 4488 10310 4502 10362
rect 4502 10310 4514 10362
rect 4514 10310 4544 10362
rect 4568 10310 4578 10362
rect 4578 10310 4624 10362
rect 4328 10308 4384 10310
rect 4408 10308 4464 10310
rect 4488 10308 4544 10310
rect 4568 10308 4624 10310
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 8758 20984 8814 21040
rect 9770 21528 9826 21584
rect 10506 21936 10562 21992
rect 10322 21528 10378 21584
rect 9678 21004 9734 21040
rect 9678 20984 9680 21004
rect 9680 20984 9732 21004
rect 9732 20984 9734 21004
rect 10138 20984 10194 21040
rect 11334 21528 11390 21584
rect 11978 22072 12034 22128
rect 12346 22072 12402 22128
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 15290 22208 15346 22264
rect 15750 21936 15806 21992
rect 14922 20848 14978 20904
rect 16486 21936 16542 21992
rect 17038 21800 17094 21856
rect 17774 22208 17830 22264
rect 19154 22228 19210 22264
rect 19154 22208 19156 22228
rect 19156 22208 19208 22228
rect 19208 22208 19210 22228
rect 20350 22108 20352 22128
rect 20352 22108 20404 22128
rect 20404 22108 20406 22128
rect 20350 22072 20406 22108
rect 18786 21836 18788 21856
rect 18788 21836 18840 21856
rect 18840 21836 18842 21856
rect 18786 21800 18842 21836
rect 9862 13812 9864 13832
rect 9864 13812 9916 13832
rect 9916 13812 9918 13832
rect 9862 13776 9918 13812
rect 10414 14220 10416 14240
rect 10416 14220 10468 14240
rect 10468 14220 10470 14240
rect 10414 14184 10470 14220
rect 11426 14184 11482 14240
rect 11058 13812 11060 13832
rect 11060 13812 11112 13832
rect 11112 13812 11114 13832
rect 11058 13776 11114 13812
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 9954 7964 9956 7984
rect 9956 7964 10008 7984
rect 10008 7964 10010 7984
rect 9954 7928 10010 7964
rect 12714 7964 12716 7984
rect 12716 7964 12768 7984
rect 12768 7964 12770 7984
rect 12714 7928 12770 7964
rect 16486 9424 16542 9480
rect 22374 22092 22430 22128
rect 22374 22072 22376 22092
rect 22376 22072 22428 22092
rect 22428 22072 22430 22092
rect 23018 19624 23074 19680
rect 20350 8880 20406 8936
rect 21362 9460 21364 9480
rect 21364 9460 21416 9480
rect 21416 9460 21418 9480
rect 21362 9424 21418 9460
rect 23018 11736 23074 11792
rect 22742 8880 22798 8936
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 22926 3848 22982 3904
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
<< metal3 >>
rect 4318 23424 4634 23425
rect 4318 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4634 23424
rect 4318 23359 4634 23360
rect 3658 22880 3974 22881
rect 3658 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3974 22880
rect 3658 22815 3974 22816
rect 4318 22336 4634 22337
rect 4318 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4634 22336
rect 4318 22271 4634 22272
rect 15285 22266 15351 22269
rect 17769 22266 17835 22269
rect 19149 22266 19215 22269
rect 15285 22264 19215 22266
rect 15285 22208 15290 22264
rect 15346 22208 17774 22264
rect 17830 22208 19154 22264
rect 19210 22208 19215 22264
rect 15285 22206 19215 22208
rect 15285 22203 15351 22206
rect 17769 22203 17835 22206
rect 19149 22203 19215 22206
rect 11973 22130 12039 22133
rect 12341 22130 12407 22133
rect 11973 22128 12407 22130
rect 11973 22072 11978 22128
rect 12034 22072 12346 22128
rect 12402 22072 12407 22128
rect 11973 22070 12407 22072
rect 11973 22067 12039 22070
rect 12341 22067 12407 22070
rect 20345 22130 20411 22133
rect 22369 22130 22435 22133
rect 20345 22128 22435 22130
rect 20345 22072 20350 22128
rect 20406 22072 22374 22128
rect 22430 22072 22435 22128
rect 20345 22070 22435 22072
rect 20345 22067 20411 22070
rect 22369 22067 22435 22070
rect 10501 21994 10567 21997
rect 15745 21994 15811 21997
rect 16481 21994 16547 21997
rect 10501 21992 16547 21994
rect 10501 21936 10506 21992
rect 10562 21936 15750 21992
rect 15806 21936 16486 21992
rect 16542 21936 16547 21992
rect 10501 21934 16547 21936
rect 10501 21931 10567 21934
rect 15745 21931 15811 21934
rect 16481 21931 16547 21934
rect 17033 21858 17099 21861
rect 18781 21858 18847 21861
rect 17033 21856 18847 21858
rect 17033 21800 17038 21856
rect 17094 21800 18786 21856
rect 18842 21800 18847 21856
rect 17033 21798 18847 21800
rect 17033 21795 17099 21798
rect 18781 21795 18847 21798
rect 3658 21792 3974 21793
rect 3658 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3974 21792
rect 3658 21727 3974 21728
rect 9765 21586 9831 21589
rect 10317 21586 10383 21589
rect 11329 21586 11395 21589
rect 9765 21584 11395 21586
rect 9765 21528 9770 21584
rect 9826 21528 10322 21584
rect 10378 21528 11334 21584
rect 11390 21528 11395 21584
rect 9765 21526 11395 21528
rect 9765 21523 9831 21526
rect 10317 21523 10383 21526
rect 11329 21523 11395 21526
rect 4318 21248 4634 21249
rect 4318 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4634 21248
rect 4318 21183 4634 21184
rect 8753 21042 8819 21045
rect 9673 21042 9739 21045
rect 10133 21042 10199 21045
rect 8753 21040 10199 21042
rect 8753 20984 8758 21040
rect 8814 20984 9678 21040
rect 9734 20984 10138 21040
rect 10194 20984 10199 21040
rect 8753 20982 10199 20984
rect 8753 20979 8819 20982
rect 9673 20979 9739 20982
rect 10133 20979 10199 20982
rect 6085 20906 6151 20909
rect 14917 20906 14983 20909
rect 6085 20904 14983 20906
rect 6085 20848 6090 20904
rect 6146 20848 14922 20904
rect 14978 20848 14983 20904
rect 6085 20846 14983 20848
rect 6085 20843 6151 20846
rect 14917 20843 14983 20846
rect 3658 20704 3974 20705
rect 3658 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3974 20704
rect 3658 20639 3974 20640
rect 4318 20160 4634 20161
rect 4318 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4634 20160
rect 4318 20095 4634 20096
rect 23013 19682 23079 19685
rect 23600 19682 24000 19712
rect 23013 19680 24000 19682
rect 23013 19624 23018 19680
rect 23074 19624 24000 19680
rect 23013 19622 24000 19624
rect 23013 19619 23079 19622
rect 3658 19616 3974 19617
rect 3658 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3974 19616
rect 23600 19592 24000 19622
rect 3658 19551 3974 19552
rect 4797 19276 4863 19277
rect 4797 19274 4844 19276
rect 4752 19272 4844 19274
rect 4908 19274 4914 19276
rect 5533 19274 5599 19277
rect 4908 19272 5599 19274
rect 4752 19216 4802 19272
rect 4908 19216 5538 19272
rect 5594 19216 5599 19272
rect 4752 19214 4844 19216
rect 4797 19212 4844 19214
rect 4908 19214 5599 19216
rect 4908 19212 4914 19214
rect 4797 19211 4863 19212
rect 5533 19211 5599 19214
rect 4318 19072 4634 19073
rect 4318 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4634 19072
rect 4318 19007 4634 19008
rect 3658 18528 3974 18529
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 4318 17984 4634 17985
rect 4318 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4634 17984
rect 4318 17919 4634 17920
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 4318 16896 4634 16897
rect 4318 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4634 16896
rect 4318 16831 4634 16832
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 4318 15808 4634 15809
rect 4318 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4634 15808
rect 4318 15743 4634 15744
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 4318 14720 4634 14721
rect 4318 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4634 14720
rect 4318 14655 4634 14656
rect 10409 14242 10475 14245
rect 11421 14242 11487 14245
rect 10409 14240 11487 14242
rect 10409 14184 10414 14240
rect 10470 14184 11426 14240
rect 11482 14184 11487 14240
rect 10409 14182 11487 14184
rect 10409 14179 10475 14182
rect 11421 14179 11487 14182
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 9857 13834 9923 13837
rect 11053 13834 11119 13837
rect 9857 13832 11119 13834
rect 9857 13776 9862 13832
rect 9918 13776 11058 13832
rect 11114 13776 11119 13832
rect 9857 13774 11119 13776
rect 9857 13771 9923 13774
rect 11053 13771 11119 13774
rect 4838 13636 4844 13700
rect 4908 13698 4914 13700
rect 5349 13698 5415 13701
rect 4908 13696 5415 13698
rect 4908 13640 5354 13696
rect 5410 13640 5415 13696
rect 4908 13638 5415 13640
rect 4908 13636 4914 13638
rect 5349 13635 5415 13638
rect 4318 13632 4634 13633
rect 4318 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4634 13632
rect 4318 13567 4634 13568
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 4318 12544 4634 12545
rect 4318 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4634 12544
rect 4318 12479 4634 12480
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 23013 11794 23079 11797
rect 23600 11794 24000 11824
rect 23013 11792 24000 11794
rect 23013 11736 23018 11792
rect 23074 11736 24000 11792
rect 23013 11734 24000 11736
rect 23013 11731 23079 11734
rect 23600 11704 24000 11734
rect 4318 11456 4634 11457
rect 4318 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4634 11456
rect 4318 11391 4634 11392
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 4318 10368 4634 10369
rect 4318 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4634 10368
rect 4318 10303 4634 10304
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 16481 9482 16547 9485
rect 21357 9482 21423 9485
rect 16481 9480 21423 9482
rect 16481 9424 16486 9480
rect 16542 9424 21362 9480
rect 21418 9424 21423 9480
rect 16481 9422 21423 9424
rect 16481 9419 16547 9422
rect 21357 9419 21423 9422
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 20345 8938 20411 8941
rect 22737 8938 22803 8941
rect 20345 8936 22803 8938
rect 20345 8880 20350 8936
rect 20406 8880 22742 8936
rect 22798 8880 22803 8936
rect 20345 8878 22803 8880
rect 20345 8875 20411 8878
rect 22737 8875 22803 8878
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 9949 7986 10015 7989
rect 12709 7986 12775 7989
rect 9949 7984 12775 7986
rect 9949 7928 9954 7984
rect 10010 7928 12714 7984
rect 12770 7928 12775 7984
rect 9949 7926 12775 7928
rect 9949 7923 10015 7926
rect 12709 7923 12775 7926
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 22921 3906 22987 3909
rect 23600 3906 24000 3936
rect 22921 3904 24000 3906
rect 22921 3848 22926 3904
rect 22982 3848 24000 3904
rect 22921 3846 24000 3848
rect 22921 3843 22987 3846
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 23600 3816 24000 3846
rect 4318 3775 4634 3776
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
<< via3 >>
rect 4324 23420 4388 23424
rect 4324 23364 4328 23420
rect 4328 23364 4384 23420
rect 4384 23364 4388 23420
rect 4324 23360 4388 23364
rect 4404 23420 4468 23424
rect 4404 23364 4408 23420
rect 4408 23364 4464 23420
rect 4464 23364 4468 23420
rect 4404 23360 4468 23364
rect 4484 23420 4548 23424
rect 4484 23364 4488 23420
rect 4488 23364 4544 23420
rect 4544 23364 4548 23420
rect 4484 23360 4548 23364
rect 4564 23420 4628 23424
rect 4564 23364 4568 23420
rect 4568 23364 4624 23420
rect 4624 23364 4628 23420
rect 4564 23360 4628 23364
rect 3664 22876 3728 22880
rect 3664 22820 3668 22876
rect 3668 22820 3724 22876
rect 3724 22820 3728 22876
rect 3664 22816 3728 22820
rect 3744 22876 3808 22880
rect 3744 22820 3748 22876
rect 3748 22820 3804 22876
rect 3804 22820 3808 22876
rect 3744 22816 3808 22820
rect 3824 22876 3888 22880
rect 3824 22820 3828 22876
rect 3828 22820 3884 22876
rect 3884 22820 3888 22876
rect 3824 22816 3888 22820
rect 3904 22876 3968 22880
rect 3904 22820 3908 22876
rect 3908 22820 3964 22876
rect 3964 22820 3968 22876
rect 3904 22816 3968 22820
rect 4324 22332 4388 22336
rect 4324 22276 4328 22332
rect 4328 22276 4384 22332
rect 4384 22276 4388 22332
rect 4324 22272 4388 22276
rect 4404 22332 4468 22336
rect 4404 22276 4408 22332
rect 4408 22276 4464 22332
rect 4464 22276 4468 22332
rect 4404 22272 4468 22276
rect 4484 22332 4548 22336
rect 4484 22276 4488 22332
rect 4488 22276 4544 22332
rect 4544 22276 4548 22332
rect 4484 22272 4548 22276
rect 4564 22332 4628 22336
rect 4564 22276 4568 22332
rect 4568 22276 4624 22332
rect 4624 22276 4628 22332
rect 4564 22272 4628 22276
rect 3664 21788 3728 21792
rect 3664 21732 3668 21788
rect 3668 21732 3724 21788
rect 3724 21732 3728 21788
rect 3664 21728 3728 21732
rect 3744 21788 3808 21792
rect 3744 21732 3748 21788
rect 3748 21732 3804 21788
rect 3804 21732 3808 21788
rect 3744 21728 3808 21732
rect 3824 21788 3888 21792
rect 3824 21732 3828 21788
rect 3828 21732 3884 21788
rect 3884 21732 3888 21788
rect 3824 21728 3888 21732
rect 3904 21788 3968 21792
rect 3904 21732 3908 21788
rect 3908 21732 3964 21788
rect 3964 21732 3968 21788
rect 3904 21728 3968 21732
rect 4324 21244 4388 21248
rect 4324 21188 4328 21244
rect 4328 21188 4384 21244
rect 4384 21188 4388 21244
rect 4324 21184 4388 21188
rect 4404 21244 4468 21248
rect 4404 21188 4408 21244
rect 4408 21188 4464 21244
rect 4464 21188 4468 21244
rect 4404 21184 4468 21188
rect 4484 21244 4548 21248
rect 4484 21188 4488 21244
rect 4488 21188 4544 21244
rect 4544 21188 4548 21244
rect 4484 21184 4548 21188
rect 4564 21244 4628 21248
rect 4564 21188 4568 21244
rect 4568 21188 4624 21244
rect 4624 21188 4628 21244
rect 4564 21184 4628 21188
rect 3664 20700 3728 20704
rect 3664 20644 3668 20700
rect 3668 20644 3724 20700
rect 3724 20644 3728 20700
rect 3664 20640 3728 20644
rect 3744 20700 3808 20704
rect 3744 20644 3748 20700
rect 3748 20644 3804 20700
rect 3804 20644 3808 20700
rect 3744 20640 3808 20644
rect 3824 20700 3888 20704
rect 3824 20644 3828 20700
rect 3828 20644 3884 20700
rect 3884 20644 3888 20700
rect 3824 20640 3888 20644
rect 3904 20700 3968 20704
rect 3904 20644 3908 20700
rect 3908 20644 3964 20700
rect 3964 20644 3968 20700
rect 3904 20640 3968 20644
rect 4324 20156 4388 20160
rect 4324 20100 4328 20156
rect 4328 20100 4384 20156
rect 4384 20100 4388 20156
rect 4324 20096 4388 20100
rect 4404 20156 4468 20160
rect 4404 20100 4408 20156
rect 4408 20100 4464 20156
rect 4464 20100 4468 20156
rect 4404 20096 4468 20100
rect 4484 20156 4548 20160
rect 4484 20100 4488 20156
rect 4488 20100 4544 20156
rect 4544 20100 4548 20156
rect 4484 20096 4548 20100
rect 4564 20156 4628 20160
rect 4564 20100 4568 20156
rect 4568 20100 4624 20156
rect 4624 20100 4628 20156
rect 4564 20096 4628 20100
rect 3664 19612 3728 19616
rect 3664 19556 3668 19612
rect 3668 19556 3724 19612
rect 3724 19556 3728 19612
rect 3664 19552 3728 19556
rect 3744 19612 3808 19616
rect 3744 19556 3748 19612
rect 3748 19556 3804 19612
rect 3804 19556 3808 19612
rect 3744 19552 3808 19556
rect 3824 19612 3888 19616
rect 3824 19556 3828 19612
rect 3828 19556 3884 19612
rect 3884 19556 3888 19612
rect 3824 19552 3888 19556
rect 3904 19612 3968 19616
rect 3904 19556 3908 19612
rect 3908 19556 3964 19612
rect 3964 19556 3968 19612
rect 3904 19552 3968 19556
rect 4844 19272 4908 19276
rect 4844 19216 4858 19272
rect 4858 19216 4908 19272
rect 4844 19212 4908 19216
rect 4324 19068 4388 19072
rect 4324 19012 4328 19068
rect 4328 19012 4384 19068
rect 4384 19012 4388 19068
rect 4324 19008 4388 19012
rect 4404 19068 4468 19072
rect 4404 19012 4408 19068
rect 4408 19012 4464 19068
rect 4464 19012 4468 19068
rect 4404 19008 4468 19012
rect 4484 19068 4548 19072
rect 4484 19012 4488 19068
rect 4488 19012 4544 19068
rect 4544 19012 4548 19068
rect 4484 19008 4548 19012
rect 4564 19068 4628 19072
rect 4564 19012 4568 19068
rect 4568 19012 4624 19068
rect 4624 19012 4628 19068
rect 4564 19008 4628 19012
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 4324 17980 4388 17984
rect 4324 17924 4328 17980
rect 4328 17924 4384 17980
rect 4384 17924 4388 17980
rect 4324 17920 4388 17924
rect 4404 17980 4468 17984
rect 4404 17924 4408 17980
rect 4408 17924 4464 17980
rect 4464 17924 4468 17980
rect 4404 17920 4468 17924
rect 4484 17980 4548 17984
rect 4484 17924 4488 17980
rect 4488 17924 4544 17980
rect 4544 17924 4548 17980
rect 4484 17920 4548 17924
rect 4564 17980 4628 17984
rect 4564 17924 4568 17980
rect 4568 17924 4624 17980
rect 4624 17924 4628 17980
rect 4564 17920 4628 17924
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 4324 16892 4388 16896
rect 4324 16836 4328 16892
rect 4328 16836 4384 16892
rect 4384 16836 4388 16892
rect 4324 16832 4388 16836
rect 4404 16892 4468 16896
rect 4404 16836 4408 16892
rect 4408 16836 4464 16892
rect 4464 16836 4468 16892
rect 4404 16832 4468 16836
rect 4484 16892 4548 16896
rect 4484 16836 4488 16892
rect 4488 16836 4544 16892
rect 4544 16836 4548 16892
rect 4484 16832 4548 16836
rect 4564 16892 4628 16896
rect 4564 16836 4568 16892
rect 4568 16836 4624 16892
rect 4624 16836 4628 16892
rect 4564 16832 4628 16836
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 4324 15804 4388 15808
rect 4324 15748 4328 15804
rect 4328 15748 4384 15804
rect 4384 15748 4388 15804
rect 4324 15744 4388 15748
rect 4404 15804 4468 15808
rect 4404 15748 4408 15804
rect 4408 15748 4464 15804
rect 4464 15748 4468 15804
rect 4404 15744 4468 15748
rect 4484 15804 4548 15808
rect 4484 15748 4488 15804
rect 4488 15748 4544 15804
rect 4544 15748 4548 15804
rect 4484 15744 4548 15748
rect 4564 15804 4628 15808
rect 4564 15748 4568 15804
rect 4568 15748 4624 15804
rect 4624 15748 4628 15804
rect 4564 15744 4628 15748
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 4324 14716 4388 14720
rect 4324 14660 4328 14716
rect 4328 14660 4384 14716
rect 4384 14660 4388 14716
rect 4324 14656 4388 14660
rect 4404 14716 4468 14720
rect 4404 14660 4408 14716
rect 4408 14660 4464 14716
rect 4464 14660 4468 14716
rect 4404 14656 4468 14660
rect 4484 14716 4548 14720
rect 4484 14660 4488 14716
rect 4488 14660 4544 14716
rect 4544 14660 4548 14716
rect 4484 14656 4548 14660
rect 4564 14716 4628 14720
rect 4564 14660 4568 14716
rect 4568 14660 4624 14716
rect 4624 14660 4628 14716
rect 4564 14656 4628 14660
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 4844 13636 4908 13700
rect 4324 13628 4388 13632
rect 4324 13572 4328 13628
rect 4328 13572 4384 13628
rect 4384 13572 4388 13628
rect 4324 13568 4388 13572
rect 4404 13628 4468 13632
rect 4404 13572 4408 13628
rect 4408 13572 4464 13628
rect 4464 13572 4468 13628
rect 4404 13568 4468 13572
rect 4484 13628 4548 13632
rect 4484 13572 4488 13628
rect 4488 13572 4544 13628
rect 4544 13572 4548 13628
rect 4484 13568 4548 13572
rect 4564 13628 4628 13632
rect 4564 13572 4568 13628
rect 4568 13572 4624 13628
rect 4624 13572 4628 13628
rect 4564 13568 4628 13572
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 4324 12540 4388 12544
rect 4324 12484 4328 12540
rect 4328 12484 4384 12540
rect 4384 12484 4388 12540
rect 4324 12480 4388 12484
rect 4404 12540 4468 12544
rect 4404 12484 4408 12540
rect 4408 12484 4464 12540
rect 4464 12484 4468 12540
rect 4404 12480 4468 12484
rect 4484 12540 4548 12544
rect 4484 12484 4488 12540
rect 4488 12484 4544 12540
rect 4544 12484 4548 12540
rect 4484 12480 4548 12484
rect 4564 12540 4628 12544
rect 4564 12484 4568 12540
rect 4568 12484 4624 12540
rect 4624 12484 4628 12540
rect 4564 12480 4628 12484
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 4324 11452 4388 11456
rect 4324 11396 4328 11452
rect 4328 11396 4384 11452
rect 4384 11396 4388 11452
rect 4324 11392 4388 11396
rect 4404 11452 4468 11456
rect 4404 11396 4408 11452
rect 4408 11396 4464 11452
rect 4464 11396 4468 11452
rect 4404 11392 4468 11396
rect 4484 11452 4548 11456
rect 4484 11396 4488 11452
rect 4488 11396 4544 11452
rect 4544 11396 4548 11452
rect 4484 11392 4548 11396
rect 4564 11452 4628 11456
rect 4564 11396 4568 11452
rect 4568 11396 4624 11452
rect 4624 11396 4628 11452
rect 4564 11392 4628 11396
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 4324 10364 4388 10368
rect 4324 10308 4328 10364
rect 4328 10308 4384 10364
rect 4384 10308 4388 10364
rect 4324 10304 4388 10308
rect 4404 10364 4468 10368
rect 4404 10308 4408 10364
rect 4408 10308 4464 10364
rect 4464 10308 4468 10364
rect 4404 10304 4468 10308
rect 4484 10364 4548 10368
rect 4484 10308 4488 10364
rect 4488 10308 4544 10364
rect 4544 10308 4548 10364
rect 4484 10304 4548 10308
rect 4564 10364 4628 10368
rect 4564 10308 4568 10364
rect 4568 10308 4624 10364
rect 4624 10308 4628 10364
rect 4564 10304 4628 10308
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
<< metal4 >>
rect 3660 23440 3980 23680
rect 3656 23420 3980 23440
rect 4316 23424 4636 23440
rect 3656 22880 3976 23420
rect 3656 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3976 22880
rect 3656 21792 3976 22816
rect 3656 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3976 21792
rect 3656 20704 3976 21728
rect 3656 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3976 20704
rect 3656 19616 3976 20640
rect 3656 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3976 19616
rect 3656 18528 3976 19552
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 3656 17440 3976 18464
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3656 15264 3976 16288
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3656 14176 3976 15200
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3656 12000 3976 13024
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4636 23424
rect 4316 22336 4636 23360
rect 4316 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4636 22336
rect 4316 21248 4636 22272
rect 4316 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4636 21248
rect 4316 20160 4636 21184
rect 4316 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4636 20160
rect 4316 19072 4636 20096
rect 4843 19276 4909 19277
rect 4843 19212 4844 19276
rect 4908 19212 4909 19276
rect 4843 19211 4909 19212
rect 4316 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4636 19072
rect 4316 17984 4636 19008
rect 4316 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4636 17984
rect 4316 16896 4636 17920
rect 4316 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4636 16896
rect 4316 15808 4636 16832
rect 4316 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4636 15808
rect 4316 14720 4636 15744
rect 4316 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4636 14720
rect 4316 13632 4636 14656
rect 4846 13701 4906 19211
rect 4843 13700 4909 13701
rect 4843 13636 4844 13700
rect 4908 13636 4909 13700
rect 4843 13635 4909 13636
rect 4316 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4636 13632
rect 4316 12544 4636 13568
rect 4316 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4636 12544
rect 4316 11456 4636 12480
rect 4316 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4636 11456
rect 4316 10368 4636 11392
rect 4316 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4636 10368
rect 4316 9280 4636 10304
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
rect 4320 320 4620 496
use sky130_fd_sc_hd__inv_2  _0490_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 23092 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1723858470
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1723858470
transform 1 0 5428 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1723858470
transform 1 0 4600 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1723858470
transform 1 0 6716 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_6  _0495_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 20424 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0496_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6072 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0497_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5888 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0498_
timestamp 1723858470
transform -1 0 9016 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0499_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9476 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0500_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 12696 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0501_
timestamp 1723858470
transform 1 0 12052 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0502_
timestamp 1723858470
transform 1 0 13892 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0503_
timestamp 1723858470
transform 1 0 14904 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0504_
timestamp 1723858470
transform 1 0 16376 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0505_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 17480 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0506_
timestamp 1723858470
transform 1 0 19136 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0507_
timestamp 1723858470
transform 1 0 20056 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0508_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21620 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0509_
timestamp 1723858470
transform 1 0 22172 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _0510_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0511_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5612 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0512_
timestamp 1723858470
transform 1 0 4048 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0513_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5060 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0514_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5060 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0515_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4600 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _0516_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4600 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0517_
timestamp 1723858470
transform 1 0 4048 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0518_
timestamp 1723858470
transform 1 0 5152 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0519_
timestamp 1723858470
transform 1 0 4876 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0520_
timestamp 1723858470
transform 1 0 4140 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0521_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4600 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0522_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5796 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0523_
timestamp 1723858470
transform 1 0 5796 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0524_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 10396 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0525_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9752 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0526_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5428 0 1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__mux2_1  _0527_
timestamp 1723858470
transform 1 0 6532 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0528_
timestamp 1723858470
transform 1 0 6440 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _0529_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4600 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0530_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5796 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0531_
timestamp 1723858470
transform 1 0 6532 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0532_
timestamp 1723858470
transform -1 0 7820 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0533_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8924 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0534_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7820 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0535_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8648 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0536_
timestamp 1723858470
transform -1 0 7452 0 1 21216
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0537_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5796 0 -1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_2  _0538_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _0539_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5428 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0540_
timestamp 1723858470
transform 1 0 7544 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0541_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6348 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0542_
timestamp 1723858470
transform 1 0 8556 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0543_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8740 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0544_
timestamp 1723858470
transform 1 0 9384 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0545_
timestamp 1723858470
transform -1 0 8740 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0546_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8280 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0547_
timestamp 1723858470
transform 1 0 7636 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0548_
timestamp 1723858470
transform -1 0 9108 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0549_
timestamp 1723858470
transform -1 0 8648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1723858470
transform -1 0 8188 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0551_
timestamp 1723858470
transform 1 0 8096 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0552_
timestamp 1723858470
transform 1 0 8188 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0553_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9936 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0554_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 12052 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0555_
timestamp 1723858470
transform -1 0 12972 0 -1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1723858470
transform -1 0 10120 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0557_
timestamp 1723858470
transform 1 0 5244 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0558_
timestamp 1723858470
transform 1 0 5796 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_2  _0559_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5244 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0560_
timestamp 1723858470
transform -1 0 7636 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0561_
timestamp 1723858470
transform 1 0 7084 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0562_
timestamp 1723858470
transform -1 0 10028 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0563_
timestamp 1723858470
transform -1 0 9384 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0564_
timestamp 1723858470
transform 1 0 9384 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0565_
timestamp 1723858470
transform -1 0 9200 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0566_
timestamp 1723858470
transform 1 0 8740 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0567_
timestamp 1723858470
transform 1 0 9200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0568_
timestamp 1723858470
transform -1 0 9384 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0569_
timestamp 1723858470
transform -1 0 9476 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0570_
timestamp 1723858470
transform 1 0 8648 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _0571_
timestamp 1723858470
transform -1 0 11316 0 1 19040
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0572_
timestamp 1723858470
transform -1 0 10856 0 -1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_1  _0573_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4692 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0574_
timestamp 1723858470
transform 1 0 5060 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0575_
timestamp 1723858470
transform 1 0 5244 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0576_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4968 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0577_
timestamp 1723858470
transform 1 0 6072 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0578_
timestamp 1723858470
transform 1 0 5796 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0579_
timestamp 1723858470
transform 1 0 7084 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0580_
timestamp 1723858470
transform 1 0 8648 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0581_
timestamp 1723858470
transform 1 0 9292 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0582_
timestamp 1723858470
transform 1 0 8648 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0583_
timestamp 1723858470
transform 1 0 9936 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0584_
timestamp 1723858470
transform -1 0 10028 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0585_
timestamp 1723858470
transform 1 0 10212 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0586_
timestamp 1723858470
transform 1 0 9568 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0587_
timestamp 1723858470
transform -1 0 10212 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0588_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9108 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0589_
timestamp 1723858470
transform 1 0 9568 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0590_
timestamp 1723858470
transform -1 0 11408 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _0591_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10948 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0592_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5428 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__o31a_1  _0593_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5152 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0594_
timestamp 1723858470
transform 1 0 4600 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0595_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5428 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0596_
timestamp 1723858470
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0597_
timestamp 1723858470
transform 1 0 5060 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0598_
timestamp 1723858470
transform 1 0 6440 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0599_
timestamp 1723858470
transform 1 0 6900 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _0600_
timestamp 1723858470
transform 1 0 6900 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0601_
timestamp 1723858470
transform 1 0 7360 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0602_
timestamp 1723858470
transform 1 0 11316 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0603_
timestamp 1723858470
transform -1 0 10856 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0604_
timestamp 1723858470
transform -1 0 10856 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0605_
timestamp 1723858470
transform -1 0 10396 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0606_
timestamp 1723858470
transform -1 0 11500 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0607_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9200 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0608_
timestamp 1723858470
transform -1 0 9384 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0609_
timestamp 1723858470
transform 1 0 10672 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _0610_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 10672 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0611_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 11500 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0612_
timestamp 1723858470
transform -1 0 11776 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0613_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10948 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0614_
timestamp 1723858470
transform -1 0 16008 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0615_
timestamp 1723858470
transform 1 0 15272 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0616_
timestamp 1723858470
transform -1 0 15640 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0617_
timestamp 1723858470
transform -1 0 16008 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0618_
timestamp 1723858470
transform 1 0 15640 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0619_
timestamp 1723858470
transform 1 0 14720 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _0620_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9016 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0621_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8924 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0622_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9200 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0623_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8280 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0624_
timestamp 1723858470
transform 1 0 10488 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0625_
timestamp 1723858470
transform 1 0 10764 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0626_
timestamp 1723858470
transform 1 0 6164 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0627_
timestamp 1723858470
transform 1 0 11776 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0628_
timestamp 1723858470
transform 1 0 11132 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0629_
timestamp 1723858470
transform 1 0 11500 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0630_
timestamp 1723858470
transform -1 0 12512 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0631_
timestamp 1723858470
transform 1 0 12512 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0632_
timestamp 1723858470
transform -1 0 12880 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0633_
timestamp 1723858470
transform -1 0 12328 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0634_
timestamp 1723858470
transform 1 0 12328 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2ai_1  _0635_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 11960 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0636_
timestamp 1723858470
transform -1 0 14536 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_4  _0637_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 16100 0 -1 22304
box -38 -48 1418 592
use sky130_fd_sc_hd__a21oi_2  _0638_
timestamp 1723858470
transform 1 0 17940 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0639_
timestamp 1723858470
transform 1 0 18676 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0640_
timestamp 1723858470
transform 1 0 19136 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0641_
timestamp 1723858470
transform 1 0 18676 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _0642_
timestamp 1723858470
transform -1 0 9844 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _0643_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9292 0 1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0644_
timestamp 1723858470
transform 1 0 12328 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0645_
timestamp 1723858470
transform -1 0 12328 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0646_
timestamp 1723858470
transform -1 0 11316 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0647_
timestamp 1723858470
transform 1 0 12788 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0648_
timestamp 1723858470
transform -1 0 12696 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0649_
timestamp 1723858470
transform 1 0 13984 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0650_
timestamp 1723858470
transform -1 0 14720 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _0651_
timestamp 1723858470
transform -1 0 12604 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0652_
timestamp 1723858470
transform 1 0 12972 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0653_
timestamp 1723858470
transform 1 0 12880 0 -1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0654_
timestamp 1723858470
transform -1 0 14260 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0655_
timestamp 1723858470
transform 1 0 13064 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0656_
timestamp 1723858470
transform 1 0 13524 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0657_
timestamp 1723858470
transform 1 0 12696 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _0658_
timestamp 1723858470
transform 1 0 18492 0 -1 22304
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_1  _0659_
timestamp 1723858470
transform 1 0 10028 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0660_
timestamp 1723858470
transform 1 0 10304 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 1723858470
transform 1 0 10488 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0662_
timestamp 1723858470
transform 1 0 7820 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0663_
timestamp 1723858470
transform 1 0 9844 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0664_
timestamp 1723858470
transform 1 0 9660 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0665_
timestamp 1723858470
transform 1 0 10948 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_1  _0666_
timestamp 1723858470
transform 1 0 12144 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0667_
timestamp 1723858470
transform 1 0 13524 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0668_
timestamp 1723858470
transform 1 0 12696 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0669_
timestamp 1723858470
transform -1 0 14628 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0670_
timestamp 1723858470
transform 1 0 13064 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0671_
timestamp 1723858470
transform -1 0 13616 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0672_
timestamp 1723858470
transform 1 0 13524 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0673_
timestamp 1723858470
transform 1 0 13616 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0674_
timestamp 1723858470
transform -1 0 13432 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0675_
timestamp 1723858470
transform 1 0 14076 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0676_
timestamp 1723858470
transform 1 0 13800 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0677_
timestamp 1723858470
transform -1 0 7912 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0678_
timestamp 1723858470
transform 1 0 8372 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0679_
timestamp 1723858470
transform 1 0 10120 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0680_
timestamp 1723858470
transform -1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0681_
timestamp 1723858470
transform 1 0 11776 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0682_
timestamp 1723858470
transform 1 0 11408 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0683_
timestamp 1723858470
transform 1 0 12512 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0684_
timestamp 1723858470
transform 1 0 12972 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0685_
timestamp 1723858470
transform -1 0 14628 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0686_
timestamp 1723858470
transform 1 0 13616 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0687_
timestamp 1723858470
transform 1 0 13524 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0688_
timestamp 1723858470
transform -1 0 14168 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0689_
timestamp 1723858470
transform -1 0 14168 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1723858470
transform 1 0 14168 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0691_
timestamp 1723858470
transform 1 0 14076 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1723858470
transform 1 0 14720 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0693_
timestamp 1723858470
transform 1 0 9476 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0694_
timestamp 1723858470
transform 1 0 7636 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0695_
timestamp 1723858470
transform 1 0 10764 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0696_
timestamp 1723858470
transform 1 0 10212 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0697_
timestamp 1723858470
transform 1 0 12144 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0698_
timestamp 1723858470
transform -1 0 13432 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0699_
timestamp 1723858470
transform 1 0 13064 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0700_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12880 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 1723858470
transform -1 0 14996 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0702_
timestamp 1723858470
transform 1 0 13524 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0703_
timestamp 1723858470
transform 1 0 14076 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1723858470
transform -1 0 16100 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0705_
timestamp 1723858470
transform 1 0 4048 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0706_
timestamp 1723858470
transform 1 0 5428 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0707_
timestamp 1723858470
transform -1 0 6348 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0708_
timestamp 1723858470
transform 1 0 5704 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0709_
timestamp 1723858470
transform 1 0 7268 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _0710_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8832 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0711_
timestamp 1723858470
transform 1 0 10672 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0712_
timestamp 1723858470
transform 1 0 10028 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0713_
timestamp 1723858470
transform 1 0 11960 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _0714_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12144 0 1 17952
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0715_
timestamp 1723858470
transform 1 0 13524 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1723858470
transform 1 0 16560 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0717_
timestamp 1723858470
transform 1 0 12788 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0718_
timestamp 1723858470
transform 1 0 14168 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0719_
timestamp 1723858470
transform -1 0 14536 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0720_
timestamp 1723858470
transform -1 0 14996 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0721_
timestamp 1723858470
transform 1 0 15180 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0722_
timestamp 1723858470
transform -1 0 15732 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0723_
timestamp 1723858470
transform -1 0 16744 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 1723858470
transform 1 0 5428 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0725_
timestamp 1723858470
transform 1 0 5428 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0726_
timestamp 1723858470
transform 1 0 5888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0727_
timestamp 1723858470
transform -1 0 5520 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0728_
timestamp 1723858470
transform 1 0 6072 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0729_
timestamp 1723858470
transform 1 0 5796 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0730_
timestamp 1723858470
transform 1 0 6992 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0731_
timestamp 1723858470
transform -1 0 7176 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0732_
timestamp 1723858470
transform 1 0 15180 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0733_
timestamp 1723858470
transform 1 0 14720 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0734_
timestamp 1723858470
transform -1 0 16008 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0735_
timestamp 1723858470
transform 1 0 11132 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0736_
timestamp 1723858470
transform -1 0 16560 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0737_
timestamp 1723858470
transform 1 0 16836 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0738_
timestamp 1723858470
transform 1 0 14812 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1723858470
transform 1 0 16560 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0740_
timestamp 1723858470
transform -1 0 17020 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0741_
timestamp 1723858470
transform -1 0 16652 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0742_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 16744 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1723858470
transform 1 0 14904 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0744_
timestamp 1723858470
transform 1 0 16284 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0745_
timestamp 1723858470
transform -1 0 16376 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0746_
timestamp 1723858470
transform 1 0 17020 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0747_
timestamp 1723858470
transform 1 0 16468 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0748_
timestamp 1723858470
transform -1 0 17204 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0749_
timestamp 1723858470
transform -1 0 7268 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0750_
timestamp 1723858470
transform 1 0 16928 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0751_
timestamp 1723858470
transform 1 0 16284 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0752_
timestamp 1723858470
transform 1 0 17204 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0753_
timestamp 1723858470
transform 1 0 16560 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0754_
timestamp 1723858470
transform -1 0 16468 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0755_
timestamp 1723858470
transform -1 0 18216 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0756_
timestamp 1723858470
transform -1 0 17940 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0757_
timestamp 1723858470
transform -1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0758_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 13708 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0759_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 16100 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _0760_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 14628 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0761_
timestamp 1723858470
transform 1 0 16100 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0762_
timestamp 1723858470
transform 1 0 16100 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0763_
timestamp 1723858470
transform 1 0 17112 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0764_
timestamp 1723858470
transform -1 0 18492 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0765_
timestamp 1723858470
transform 1 0 18308 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0766_
timestamp 1723858470
transform 1 0 18768 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _0767_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 18032 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0768_
timestamp 1723858470
transform -1 0 18124 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0769_
timestamp 1723858470
transform -1 0 17572 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0770_
timestamp 1723858470
transform 1 0 17480 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0771_
timestamp 1723858470
transform 1 0 17664 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1723858470
transform 1 0 18676 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0773_
timestamp 1723858470
transform -1 0 18216 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0774_
timestamp 1723858470
transform 1 0 17572 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0775_
timestamp 1723858470
transform -1 0 18216 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0776_
timestamp 1723858470
transform -1 0 18492 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0777_
timestamp 1723858470
transform 1 0 17664 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0778_
timestamp 1723858470
transform -1 0 19320 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0779_
timestamp 1723858470
transform 1 0 19320 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0780_
timestamp 1723858470
transform 1 0 20516 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0781_
timestamp 1723858470
transform -1 0 20516 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0782_
timestamp 1723858470
transform 1 0 20608 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0783_
timestamp 1723858470
transform 1 0 21252 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0784_
timestamp 1723858470
transform 1 0 21712 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0785_
timestamp 1723858470
transform -1 0 21804 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0786_
timestamp 1723858470
transform 1 0 20976 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0787_
timestamp 1723858470
transform 1 0 18216 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _0788_
timestamp 1723858470
transform 1 0 20516 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0789_
timestamp 1723858470
transform -1 0 20516 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1723858470
transform 1 0 20056 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o311ai_2  _0791_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 17112 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0792_
timestamp 1723858470
transform 1 0 18676 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0793_
timestamp 1723858470
transform -1 0 18676 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0794_
timestamp 1723858470
transform -1 0 19504 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0795_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0796_
timestamp 1723858470
transform -1 0 20424 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0797_
timestamp 1723858470
transform 1 0 19504 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0798_
timestamp 1723858470
transform -1 0 22724 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0799_
timestamp 1723858470
transform -1 0 20424 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0800_
timestamp 1723858470
transform 1 0 21804 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _0801_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21160 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0802_
timestamp 1723858470
transform -1 0 21804 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0803_
timestamp 1723858470
transform -1 0 20700 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0804_
timestamp 1723858470
transform -1 0 21160 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0805_
timestamp 1723858470
transform 1 0 20516 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0806_
timestamp 1723858470
transform -1 0 21160 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0807_
timestamp 1723858470
transform 1 0 21252 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0808_
timestamp 1723858470
transform 1 0 20976 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0809_
timestamp 1723858470
transform -1 0 21068 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0810_
timestamp 1723858470
transform -1 0 22908 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0811_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21252 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0812_
timestamp 1723858470
transform 1 0 19964 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0813_
timestamp 1723858470
transform -1 0 22816 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0814_
timestamp 1723858470
transform 1 0 21528 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0815_
timestamp 1723858470
transform 1 0 21620 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0816_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 20516 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0817_
timestamp 1723858470
transform 1 0 21252 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0818_
timestamp 1723858470
transform -1 0 21620 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0819_
timestamp 1723858470
transform 1 0 21528 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0820_
timestamp 1723858470
transform 1 0 20976 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0821_
timestamp 1723858470
transform 1 0 21160 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0822_
timestamp 1723858470
transform 1 0 20516 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0823_
timestamp 1723858470
transform 1 0 20240 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0824_
timestamp 1723858470
transform -1 0 21068 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0825_
timestamp 1723858470
transform -1 0 19964 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1723858470
transform -1 0 19780 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0827_
timestamp 1723858470
transform 1 0 19412 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0828_
timestamp 1723858470
transform -1 0 19320 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0829_
timestamp 1723858470
transform 1 0 18308 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0830_
timestamp 1723858470
transform -1 0 17848 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0831_
timestamp 1723858470
transform 1 0 17848 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0832_
timestamp 1723858470
transform -1 0 18308 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0833_
timestamp 1723858470
transform 1 0 18676 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0834_
timestamp 1723858470
transform 1 0 16836 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0835_
timestamp 1723858470
transform 1 0 17204 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0836_
timestamp 1723858470
transform -1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1723858470
transform 1 0 17756 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0838_
timestamp 1723858470
transform 1 0 16100 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0839_
timestamp 1723858470
transform 1 0 16376 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0840_
timestamp 1723858470
transform 1 0 14628 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0841_
timestamp 1723858470
transform -1 0 17480 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0842_
timestamp 1723858470
transform -1 0 16560 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0843_
timestamp 1723858470
transform 1 0 14076 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0844_
timestamp 1723858470
transform 1 0 14812 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0845_
timestamp 1723858470
transform 1 0 14168 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0846_
timestamp 1723858470
transform 1 0 14720 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0847_
timestamp 1723858470
transform 1 0 14168 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0848_
timestamp 1723858470
transform 1 0 11500 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0849_
timestamp 1723858470
transform 1 0 13064 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0850_
timestamp 1723858470
transform 1 0 13524 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0851_
timestamp 1723858470
transform 1 0 11224 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0852_
timestamp 1723858470
transform 1 0 11592 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0853_
timestamp 1723858470
transform 1 0 11868 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0854_
timestamp 1723858470
transform 1 0 12328 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0855_
timestamp 1723858470
transform 1 0 11132 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0856_
timestamp 1723858470
transform 1 0 9200 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0857_
timestamp 1723858470
transform 1 0 10948 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0858_
timestamp 1723858470
transform 1 0 8188 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0859_
timestamp 1723858470
transform -1 0 9476 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0860_
timestamp 1723858470
transform -1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0861_
timestamp 1723858470
transform -1 0 9016 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0862_
timestamp 1723858470
transform 1 0 8188 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0863_
timestamp 1723858470
transform 1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0864_
timestamp 1723858470
transform 1 0 7084 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0865_
timestamp 1723858470
transform -1 0 7912 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0866_
timestamp 1723858470
transform -1 0 5796 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0867_
timestamp 1723858470
transform 1 0 5152 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0868_
timestamp 1723858470
transform -1 0 7176 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0869_
timestamp 1723858470
transform 1 0 4876 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0870_
timestamp 1723858470
transform 1 0 5796 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0871_
timestamp 1723858470
transform -1 0 3680 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0872_
timestamp 1723858470
transform -1 0 3772 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0873_
timestamp 1723858470
transform 1 0 5796 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1723858470
transform 1 0 5428 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 1723858470
transform 1 0 5336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0876_
timestamp 1723858470
transform -1 0 6348 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0877_
timestamp 1723858470
transform 1 0 6072 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0878_
timestamp 1723858470
transform 1 0 7268 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0879_
timestamp 1723858470
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0880_
timestamp 1723858470
transform 1 0 12236 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0881_
timestamp 1723858470
transform 1 0 15456 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0882_
timestamp 1723858470
transform 1 0 16560 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0883_
timestamp 1723858470
transform 1 0 18952 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0884_
timestamp 1723858470
transform 1 0 20240 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0885_
timestamp 1723858470
transform -1 0 22356 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0886_
timestamp 1723858470
transform -1 0 22724 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0887_
timestamp 1723858470
transform 1 0 22356 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0888_
timestamp 1723858470
transform -1 0 22264 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0889_
timestamp 1723858470
transform 1 0 3036 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0890_
timestamp 1723858470
transform -1 0 6072 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0891_
timestamp 1723858470
transform 1 0 4692 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1723858470
transform 1 0 3772 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0893_
timestamp 1723858470
transform 1 0 3680 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0894_
timestamp 1723858470
transform -1 0 4232 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0895_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4692 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0896_
timestamp 1723858470
transform 1 0 3220 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0897_
timestamp 1723858470
transform 1 0 3496 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0898_
timestamp 1723858470
transform -1 0 4140 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0899_
timestamp 1723858470
transform -1 0 6808 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0900_
timestamp 1723858470
transform 1 0 4784 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0901_
timestamp 1723858470
transform -1 0 4784 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0902_
timestamp 1723858470
transform 1 0 5060 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0903_
timestamp 1723858470
transform -1 0 6624 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0904_
timestamp 1723858470
transform 1 0 5520 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0905_
timestamp 1723858470
transform 1 0 6716 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0906_
timestamp 1723858470
transform -1 0 7452 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0907_
timestamp 1723858470
transform 1 0 6348 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0908_
timestamp 1723858470
transform 1 0 6992 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 1723858470
transform 1 0 7728 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0910_
timestamp 1723858470
transform 1 0 7452 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0911_
timestamp 1723858470
transform 1 0 8096 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1723858470
transform 1 0 8372 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0913_
timestamp 1723858470
transform -1 0 9384 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0914_
timestamp 1723858470
transform -1 0 11224 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1723858470
transform -1 0 10856 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0916_
timestamp 1723858470
transform 1 0 9844 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0917_
timestamp 1723858470
transform -1 0 11316 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0918_
timestamp 1723858470
transform 1 0 10304 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0919_
timestamp 1723858470
transform -1 0 10856 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0920_
timestamp 1723858470
transform 1 0 11224 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0921_
timestamp 1723858470
transform 1 0 11408 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0922_
timestamp 1723858470
transform 1 0 11868 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1723858470
transform -1 0 13432 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0924_
timestamp 1723858470
transform -1 0 13800 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0925_
timestamp 1723858470
transform 1 0 12972 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0926_
timestamp 1723858470
transform 1 0 14352 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0927_
timestamp 1723858470
transform -1 0 13524 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0928_
timestamp 1723858470
transform -1 0 14352 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0929_
timestamp 1723858470
transform 1 0 14444 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0930_
timestamp 1723858470
transform 1 0 14996 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0931_
timestamp 1723858470
transform -1 0 15640 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0932_
timestamp 1723858470
transform -1 0 18124 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0933_
timestamp 1723858470
transform 1 0 16468 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0934_
timestamp 1723858470
transform -1 0 17388 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0935_
timestamp 1723858470
transform -1 0 17848 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0936_
timestamp 1723858470
transform -1 0 16652 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0937_
timestamp 1723858470
transform -1 0 17388 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0938_
timestamp 1723858470
transform -1 0 17848 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0939_
timestamp 1723858470
transform 1 0 17848 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0940_
timestamp 1723858470
transform 1 0 17480 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0941_
timestamp 1723858470
transform 1 0 16928 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0942_
timestamp 1723858470
transform -1 0 18308 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0943_
timestamp 1723858470
transform 1 0 17204 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1723858470
transform 1 0 18216 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0945_
timestamp 1723858470
transform 1 0 18676 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0946_
timestamp 1723858470
transform -1 0 18492 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0947_
timestamp 1723858470
transform 1 0 20608 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1723858470
transform -1 0 20148 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0949_
timestamp 1723858470
transform -1 0 20240 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0950_
timestamp 1723858470
transform -1 0 20884 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0951_
timestamp 1723858470
transform -1 0 20608 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0952_
timestamp 1723858470
transform -1 0 20240 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0953_
timestamp 1723858470
transform 1 0 21528 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0954_
timestamp 1723858470
transform -1 0 20884 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0955_
timestamp 1723858470
transform -1 0 21528 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0956_
timestamp 1723858470
transform 1 0 21988 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0957_
timestamp 1723858470
transform 1 0 21528 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0958_
timestamp 1723858470
transform 1 0 21436 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0959_
timestamp 1723858470
transform -1 0 22540 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0960_
timestamp 1723858470
transform 1 0 22448 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0961_
timestamp 1723858470
transform 1 0 20884 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0962_
timestamp 1723858470
transform 1 0 20332 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0963_
timestamp 1723858470
transform -1 0 22356 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0964_
timestamp 1723858470
transform 1 0 20792 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0965_
timestamp 1723858470
transform 1 0 20700 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0966_
timestamp 1723858470
transform -1 0 21804 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0967_
timestamp 1723858470
transform -1 0 21804 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0968_
timestamp 1723858470
transform -1 0 21160 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0969_
timestamp 1723858470
transform -1 0 21712 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0970_
timestamp 1723858470
transform 1 0 21804 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0971_
timestamp 1723858470
transform -1 0 22816 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0972_
timestamp 1723858470
transform -1 0 20792 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1723858470
transform -1 0 18584 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0974_
timestamp 1723858470
transform -1 0 19688 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0975_
timestamp 1723858470
transform -1 0 19412 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0976_
timestamp 1723858470
transform -1 0 19688 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0977_
timestamp 1723858470
transform 1 0 19412 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1723858470
transform -1 0 19228 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0979_
timestamp 1723858470
transform -1 0 23092 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0980_
timestamp 1723858470
transform -1 0 21620 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0981_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5612 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1723858470
transform 1 0 4232 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1723858470
transform 1 0 4232 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1723858470
transform 1 0 4508 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1723858470
transform 1 0 5980 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1723858470
transform 1 0 8372 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1723858470
transform 1 0 8096 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1723858470
transform 1 0 10948 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1723858470
transform 1 0 10672 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1723858470
transform 1 0 11776 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1723858470
transform 1 0 13524 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1723858470
transform 1 0 13432 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1723858470
transform 1 0 14352 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1723858470
transform -1 0 16008 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1723858470
transform 1 0 15640 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1723858470
transform 1 0 16100 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1723858470
transform 1 0 18676 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1723858470
transform -1 0 20056 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1723858470
transform 1 0 19136 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1723858470
transform 1 0 21252 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1723858470
transform 1 0 21344 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1723858470
transform 1 0 20792 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1723858470
transform 1 0 3864 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1723858470
transform -1 0 5796 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1723858470
transform 1 0 4232 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1723858470
transform 1 0 4140 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1723858470
transform 1 0 3588 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1723858470
transform 1 0 3956 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1723858470
transform 1 0 5796 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1723858470
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1723858470
transform -1 0 9016 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1723858470
transform 1 0 8372 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1723858470
transform 1 0 10948 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1723858470
transform 1 0 9844 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1723858470
transform -1 0 12788 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1723858470
transform 1 0 13524 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1723858470
transform -1 0 14996 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1723858470
transform -1 0 16376 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1723858470
transform 1 0 16376 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1723858470
transform -1 0 18124 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1723858470
transform -1 0 18584 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1723858470
transform 1 0 19136 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1723858470
transform 1 0 17664 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1723858470
transform 1 0 19412 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1723858470
transform 1 0 19412 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1723858470
transform 1 0 20332 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1723858470
transform -1 0 23092 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1723858470
transform 1 0 21528 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1723858470
transform 1 0 21436 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1723858470
transform 1 0 21252 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1723858470
transform 1 0 21252 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1723858470
transform 1 0 19688 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1723858470
transform 1 0 18676 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1723858470
transform 1 0 18492 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1723858470
transform 1 0 21620 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  fanout11 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12880 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout12
timestamp 1723858470
transform -1 0 22908 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout13
timestamp 1723858470
transform 1 0 21252 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout14 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21988 0 1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout15 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 20148 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout16 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 21712 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout17 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 17020 0 1 22304
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp 1723858470
transform -1 0 5520 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 1723858470
transform -1 0 4508 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1723858470
transform -1 0 5152 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1723858470
transform -1 0 21160 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1723858470
transform -1 0 22816 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout23
timestamp 1723858470
transform -1 0 9200 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout24 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8096 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1723858470
transform -1 0 12236 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1723858470
transform -1 0 23092 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1723858470
transform -1 0 16652 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1723858470
transform -1 0 22632 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp 1723858470
transform -1 0 22080 0 1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1723858470
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1723858470
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1723858470
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1723858470
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1723858470
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1723858470
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1723858470
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1723858470
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1723858470
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1723858470
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1723858470
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1723858470
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1723858470
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1723858470
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1723858470
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1723858470
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1723858470
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1723858470
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1723858470
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1723858470
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1723858470
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1723858470
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_237 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 22356 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1723858470
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1723858470
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1723858470
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1723858470
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1723858470
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1723858470
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1723858470
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1723858470
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1723858470
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1723858470
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1723858470
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1723858470
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1723858470
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1723858470
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1723858470
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1723858470
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1723858470
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1723858470
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1723858470
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1723858470
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1723858470
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1723858470
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1723858470
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_237
timestamp 1723858470
transform 1 0 22356 0 -1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1723858470
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1723858470
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1723858470
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1723858470
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1723858470
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1723858470
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1723858470
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1723858470
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1723858470
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1723858470
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1723858470
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1723858470
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1723858470
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1723858470
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1723858470
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1723858470
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1723858470
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1723858470
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1723858470
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1723858470
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1723858470
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1723858470
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1723858470
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1723858470
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1723858470
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1723858470
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1723858470
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1723858470
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1723858470
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1723858470
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1723858470
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1723858470
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1723858470
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1723858470
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1723858470
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1723858470
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1723858470
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1723858470
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1723858470
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1723858470
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1723858470
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1723858470
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1723858470
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1723858470
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1723858470
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1723858470
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1723858470
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1723858470
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1723858470
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1723858470
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_237
timestamp 1723858470
transform 1 0 22356 0 -1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1723858470
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1723858470
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1723858470
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1723858470
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1723858470
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1723858470
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1723858470
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1723858470
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1723858470
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1723858470
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1723858470
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1723858470
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1723858470
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1723858470
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1723858470
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1723858470
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1723858470
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1723858470
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1723858470
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1723858470
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1723858470
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1723858470
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1723858470
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1723858470
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1723858470
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1723858470
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1723858470
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1723858470
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1723858470
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1723858470
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1723858470
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1723858470
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1723858470
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1723858470
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1723858470
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1723858470
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1723858470
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1723858470
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1723858470
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1723858470
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1723858470
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1723858470
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1723858470
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1723858470
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1723858470
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1723858470
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1723858470
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1723858470
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1723858470
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1723858470
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_237
timestamp 1723858470
transform 1 0 22356 0 -1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1723858470
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1723858470
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1723858470
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1723858470
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1723858470
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1723858470
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1723858470
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1723858470
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1723858470
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1723858470
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1723858470
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1723858470
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1723858470
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1723858470
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1723858470
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1723858470
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1723858470
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1723858470
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1723858470
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1723858470
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1723858470
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1723858470
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1723858470
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1723858470
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_233
timestamp 1723858470
transform 1 0 21988 0 1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1723858470
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1723858470
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1723858470
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1723858470
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1723858470
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1723858470
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1723858470
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1723858470
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1723858470
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1723858470
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1723858470
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1723858470
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1723858470
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1723858470
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1723858470
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1723858470
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1723858470
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1723858470
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1723858470
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1723858470
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1723858470
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1723858470
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1723858470
transform 1 0 20516 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1723858470
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1723858470
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_237
timestamp 1723858470
transform 1 0 22356 0 -1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1723858470
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1723858470
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1723858470
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1723858470
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1723858470
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1723858470
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1723858470
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1723858470
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1723858470
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1723858470
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1723858470
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1723858470
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1723858470
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1723858470
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1723858470
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1723858470
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1723858470
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1723858470
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1723858470
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1723858470
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1723858470
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1723858470
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1723858470
transform 1 0 19780 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1723858470
transform 1 0 20884 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1723858470
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1723858470
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1723858470
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_27
timestamp 1723858470
transform 1 0 3036 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_35
timestamp 1723858470
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_52
timestamp 1723858470
transform 1 0 5336 0 -1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1723858470
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1723858470
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1723858470
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1723858470
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1723858470
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1723858470
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1723858470
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1723858470
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1723858470
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1723858470
transform 1 0 14260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1723858470
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1723858470
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1723858470
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1723858470
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1723858470
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1723858470
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1723858470
transform 1 0 20516 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1723858470
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1723858470
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_237
timestamp 1723858470
transform 1 0 22356 0 -1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1723858470
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1723858470
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1723858470
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_57
timestamp 1723858470
transform 1 0 5796 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_69
timestamp 1723858470
transform 1 0 6900 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1723858470
transform 1 0 8004 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1723858470
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_97
timestamp 1723858470
transform 1 0 9476 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_105
timestamp 1723858470
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_112
timestamp 1723858470
transform 1 0 10856 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_124
timestamp 1723858470
transform 1 0 11960 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_136
timestamp 1723858470
transform 1 0 13064 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1723858470
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1723858470
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1723858470
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1723858470
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1723858470
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1723858470
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1723858470
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1723858470
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1723858470
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1723858470
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1723858470
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1723858470
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_64
timestamp 1723858470
transform 1 0 6440 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_75
timestamp 1723858470
transform 1 0 7452 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_92
timestamp 1723858470
transform 1 0 9016 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_104
timestamp 1723858470
transform 1 0 10120 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_129
timestamp 1723858470
transform 1 0 12420 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_137
timestamp 1723858470
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_144
timestamp 1723858470
transform 1 0 13800 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_156
timestamp 1723858470
transform 1 0 14904 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1723858470
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1723858470
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1723858470
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1723858470
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1723858470
transform 1 0 20516 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1723858470
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1723858470
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_237
timestamp 1723858470
transform 1 0 22356 0 -1 7072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1723858470
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1723858470
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1723858470
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1723858470
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_60
timestamp 1723858470
transform 1 0 6072 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_133
timestamp 1723858470
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_162
timestamp 1723858470
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_174
timestamp 1723858470
transform 1 0 16560 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_186
timestamp 1723858470
transform 1 0 17664 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_194
timestamp 1723858470
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_197
timestamp 1723858470
transform 1 0 18676 0 1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_208
timestamp 1723858470
transform 1 0 19688 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_220
timestamp 1723858470
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_234
timestamp 1723858470
transform 1 0 22080 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_242
timestamp 1723858470
transform 1 0 22816 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1723858470
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1723858470
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_27
timestamp 1723858470
transform 1 0 3036 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_35
timestamp 1723858470
transform 1 0 3772 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_50
timestamp 1723858470
transform 1 0 5152 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1723858470
transform 1 0 5796 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 1723858470
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_96
timestamp 1723858470
transform 1 0 9384 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_100
timestamp 1723858470
transform 1 0 9752 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_134
timestamp 1723858470
transform 1 0 12880 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_164
timestamp 1723858470
transform 1 0 15640 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_169
timestamp 1723858470
transform 1 0 16100 0 -1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_183
timestamp 1723858470
transform 1 0 17388 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_195
timestamp 1723858470
transform 1 0 18492 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1723858470
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1723858470
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1723858470
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1723858470
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1723858470
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_53
timestamp 1723858470
transform 1 0 5428 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_66
timestamp 1723858470
transform 1 0 6624 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_94
timestamp 1723858470
transform 1 0 9200 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_106
timestamp 1723858470
transform 1 0 10304 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_117
timestamp 1723858470
transform 1 0 11316 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_127
timestamp 1723858470
transform 1 0 12236 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_135
timestamp 1723858470
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1723858470
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_155
timestamp 1723858470
transform 1 0 14812 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_220
timestamp 1723858470
transform 1 0 20792 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_242
timestamp 1723858470
transform 1 0 22816 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1723858470
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1723858470
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_27
timestamp 1723858470
transform 1 0 3036 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_73
timestamp 1723858470
transform 1 0 7268 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_81
timestamp 1723858470
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_90
timestamp 1723858470
transform 1 0 8832 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_97
timestamp 1723858470
transform 1 0 9476 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1723858470
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_133
timestamp 1723858470
transform 1 0 12788 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_145
timestamp 1723858470
transform 1 0 13892 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_158
timestamp 1723858470
transform 1 0 15088 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp 1723858470
transform 1 0 15824 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1723858470
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_175
timestamp 1723858470
transform 1 0 16652 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_188
timestamp 1723858470
transform 1 0 17848 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_194
timestamp 1723858470
transform 1 0 18400 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_241
timestamp 1723858470
transform 1 0 22724 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1723858470
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1723858470
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1723858470
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_68
timestamp 1723858470
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_72
timestamp 1723858470
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_78
timestamp 1723858470
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_92
timestamp 1723858470
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_101
timestamp 1723858470
transform 1 0 9844 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_113
timestamp 1723858470
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_122
timestamp 1723858470
transform 1 0 11776 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_134
timestamp 1723858470
transform 1 0 12880 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_168
timestamp 1723858470
transform 1 0 16008 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_191
timestamp 1723858470
transform 1 0 18124 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1723858470
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_197
timestamp 1723858470
transform 1 0 18676 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_208
timestamp 1723858470
transform 1 0 19688 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_214
timestamp 1723858470
transform 1 0 20240 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_243
timestamp 1723858470
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1723858470
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1723858470
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_27
timestamp 1723858470
transform 1 0 3036 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_33
timestamp 1723858470
transform 1 0 3588 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1723858470
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_64
timestamp 1723858470
transform 1 0 6440 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_70
timestamp 1723858470
transform 1 0 6992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_80
timestamp 1723858470
transform 1 0 7912 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_97
timestamp 1723858470
transform 1 0 9476 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1723858470
transform 1 0 10580 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_113
timestamp 1723858470
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_131
timestamp 1723858470
transform 1 0 12604 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_143
timestamp 1723858470
transform 1 0 13708 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_157
timestamp 1723858470
transform 1 0 14996 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 1723858470
transform 1 0 15732 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1723858470
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1723858470
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1723858470
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_217
timestamp 1723858470
transform 1 0 20516 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_242
timestamp 1723858470
transform 1 0 22816 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1723858470
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1723858470
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1723858470
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1723858470
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_41
timestamp 1723858470
transform 1 0 4324 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_49
timestamp 1723858470
transform 1 0 5060 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_75
timestamp 1723858470
transform 1 0 7452 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1723858470
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 1723858470
transform 1 0 8372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_103
timestamp 1723858470
transform 1 0 10028 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_118
timestamp 1723858470
transform 1 0 11408 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_135
timestamp 1723858470
transform 1 0 12972 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1723858470
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_141
timestamp 1723858470
transform 1 0 13524 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_159
timestamp 1723858470
transform 1 0 15180 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_167
timestamp 1723858470
transform 1 0 15916 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1723858470
transform 1 0 18676 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_214
timestamp 1723858470
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_231
timestamp 1723858470
transform 1 0 21804 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_239
timestamp 1723858470
transform 1 0 22540 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1723858470
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1723858470
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1723858470
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_39
timestamp 1723858470
transform 1 0 4140 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1723858470
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_57
timestamp 1723858470
transform 1 0 5796 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_65
timestamp 1723858470
transform 1 0 6532 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_77
timestamp 1723858470
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_98
timestamp 1723858470
transform 1 0 9568 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 1723858470
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_129
timestamp 1723858470
transform 1 0 12420 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_137
timestamp 1723858470
transform 1 0 13156 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_163
timestamp 1723858470
transform 1 0 15548 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1723858470
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1723858470
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_191
timestamp 1723858470
transform 1 0 18124 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_203
timestamp 1723858470
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_221
timestamp 1723858470
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_225
timestamp 1723858470
transform 1 0 21252 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_243
timestamp 1723858470
transform 1 0 22908 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1723858470
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1723858470
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1723858470
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1723858470
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1723858470
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_57
timestamp 1723858470
transform 1 0 5796 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_69
timestamp 1723858470
transform 1 0 6900 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 1723858470
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_101
timestamp 1723858470
transform 1 0 9844 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_109
timestamp 1723858470
transform 1 0 10580 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_126
timestamp 1723858470
transform 1 0 12144 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1723858470
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_141
timestamp 1723858470
transform 1 0 13524 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_166
timestamp 1723858470
transform 1 0 15824 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_178
timestamp 1723858470
transform 1 0 16928 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_186
timestamp 1723858470
transform 1 0 17664 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_193
timestamp 1723858470
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_197
timestamp 1723858470
transform 1 0 18676 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_205
timestamp 1723858470
transform 1 0 19412 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_244
timestamp 1723858470
transform 1 0 23000 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1723858470
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1723858470
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1723858470
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_39
timestamp 1723858470
transform 1 0 4140 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_57
timestamp 1723858470
transform 1 0 5796 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_63
timestamp 1723858470
transform 1 0 6348 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_73
timestamp 1723858470
transform 1 0 7268 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_79
timestamp 1723858470
transform 1 0 7820 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_97
timestamp 1723858470
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1723858470
transform 1 0 10212 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1723858470
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 1723858470
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_138
timestamp 1723858470
transform 1 0 13248 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_146
timestamp 1723858470
transform 1 0 13984 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_152
timestamp 1723858470
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_163
timestamp 1723858470
transform 1 0 15548 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1723858470
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_176
timestamp 1723858470
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1723858470
transform 1 0 21068 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1723858470
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1723858470
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1723858470
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1723858470
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_41
timestamp 1723858470
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_75
timestamp 1723858470
transform 1 0 7452 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1723858470
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1723858470
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_96
timestamp 1723858470
transform 1 0 9384 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_108
timestamp 1723858470
transform 1 0 10488 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_112
timestamp 1723858470
transform 1 0 10856 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_120
timestamp 1723858470
transform 1 0 11592 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_131
timestamp 1723858470
transform 1 0 12604 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1723858470
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_157
timestamp 1723858470
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_169
timestamp 1723858470
transform 1 0 16100 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_181
timestamp 1723858470
transform 1 0 17204 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_187
timestamp 1723858470
transform 1 0 17756 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1723858470
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_203
timestamp 1723858470
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_243
timestamp 1723858470
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1723858470
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1723858470
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1723858470
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_39
timestamp 1723858470
transform 1 0 4140 0 -1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_66
timestamp 1723858470
transform 1 0 6624 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_78
timestamp 1723858470
transform 1 0 7728 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_86
timestamp 1723858470
transform 1 0 8464 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_97
timestamp 1723858470
transform 1 0 9476 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_108
timestamp 1723858470
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1723858470
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_125
timestamp 1723858470
transform 1 0 12052 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_134
timestamp 1723858470
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_148
timestamp 1723858470
transform 1 0 14168 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_169
timestamp 1723858470
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_181
timestamp 1723858470
transform 1 0 17204 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_197
timestamp 1723858470
transform 1 0 18676 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_205
timestamp 1723858470
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_221
timestamp 1723858470
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_225
timestamp 1723858470
transform 1 0 21252 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_243
timestamp 1723858470
transform 1 0 22908 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1723858470
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1723858470
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1723858470
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1723858470
transform 1 0 3220 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_37
timestamp 1723858470
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_64
timestamp 1723858470
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_76
timestamp 1723858470
transform 1 0 7544 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_88
timestamp 1723858470
transform 1 0 8648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_119
timestamp 1723858470
transform 1 0 11500 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_135
timestamp 1723858470
transform 1 0 12972 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1723858470
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_151
timestamp 1723858470
transform 1 0 14444 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_159
timestamp 1723858470
transform 1 0 15180 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_169
timestamp 1723858470
transform 1 0 16100 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_190
timestamp 1723858470
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_202
timestamp 1723858470
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_214
timestamp 1723858470
transform 1 0 20240 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_236
timestamp 1723858470
transform 1 0 22264 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_244
timestamp 1723858470
transform 1 0 23000 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1723858470
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1723858470
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1723858470
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_39
timestamp 1723858470
transform 1 0 4140 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1723858470
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_69
timestamp 1723858470
transform 1 0 6900 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_89
timestamp 1723858470
transform 1 0 8740 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_96
timestamp 1723858470
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_119
timestamp 1723858470
transform 1 0 11500 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_131
timestamp 1723858470
transform 1 0 12604 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1723858470
transform 1 0 14260 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1723858470
transform 1 0 15364 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1723858470
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_206
timestamp 1723858470
transform 1 0 19504 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_218
timestamp 1723858470
transform 1 0 20608 0 -1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1723858470
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1723858470
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1723858470
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1723858470
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_41
timestamp 1723858470
transform 1 0 4324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_53
timestamp 1723858470
transform 1 0 5428 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_59
timestamp 1723858470
transform 1 0 5980 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_66
timestamp 1723858470
transform 1 0 6624 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 1723858470
transform 1 0 8004 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 1723858470
transform 1 0 8372 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_93
timestamp 1723858470
transform 1 0 9108 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_103
timestamp 1723858470
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_112
timestamp 1723858470
transform 1 0 10856 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_116
timestamp 1723858470
transform 1 0 11224 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_120
timestamp 1723858470
transform 1 0 11592 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_135
timestamp 1723858470
transform 1 0 12972 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1723858470
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_148
timestamp 1723858470
transform 1 0 14168 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_160
timestamp 1723858470
transform 1 0 15272 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_180
timestamp 1723858470
transform 1 0 17112 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1723858470
transform 1 0 18308 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_204
timestamp 1723858470
transform 1 0 19320 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_212
timestamp 1723858470
transform 1 0 20056 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_220
timestamp 1723858470
transform 1 0 20792 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_241
timestamp 1723858470
transform 1 0 22724 0 1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1723858470
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1723858470
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_27
timestamp 1723858470
transform 1 0 3036 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_35
timestamp 1723858470
transform 1 0 3772 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_43
timestamp 1723858470
transform 1 0 4508 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_78
timestamp 1723858470
transform 1 0 7728 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_86
timestamp 1723858470
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_100
timestamp 1723858470
transform 1 0 9752 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_107
timestamp 1723858470
transform 1 0 10396 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1723858470
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_113
timestamp 1723858470
transform 1 0 10948 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_126
timestamp 1723858470
transform 1 0 12144 0 -1 15776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_147
timestamp 1723858470
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_159
timestamp 1723858470
transform 1 0 15180 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1723858470
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_183
timestamp 1723858470
transform 1 0 17388 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_195
timestamp 1723858470
transform 1 0 18492 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_203
timestamp 1723858470
transform 1 0 19228 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_209
timestamp 1723858470
transform 1 0 19780 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_213
timestamp 1723858470
transform 1 0 20148 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1723858470
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_225
timestamp 1723858470
transform 1 0 21252 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_235
timestamp 1723858470
transform 1 0 22172 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_243
timestamp 1723858470
transform 1 0 22908 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1723858470
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1723858470
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1723858470
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1723858470
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_41
timestamp 1723858470
transform 1 0 4324 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_59
timestamp 1723858470
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_73
timestamp 1723858470
transform 1 0 7268 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 1723858470
transform 1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1723858470
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1723858470
transform 1 0 9476 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_109
timestamp 1723858470
transform 1 0 10580 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_131
timestamp 1723858470
transform 1 0 12604 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_152
timestamp 1723858470
transform 1 0 14536 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_165
timestamp 1723858470
transform 1 0 15732 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_179
timestamp 1723858470
transform 1 0 17020 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_191
timestamp 1723858470
transform 1 0 18124 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1723858470
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 1723858470
transform 1 0 18676 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_201
timestamp 1723858470
transform 1 0 19044 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_211
timestamp 1723858470
transform 1 0 19964 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_220
timestamp 1723858470
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_240
timestamp 1723858470
transform 1 0 22632 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_244
timestamp 1723858470
transform 1 0 23000 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1723858470
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1723858470
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1723858470
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1723858470
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_69
timestamp 1723858470
transform 1 0 6900 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_80
timestamp 1723858470
transform 1 0 7912 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_88
timestamp 1723858470
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_101
timestamp 1723858470
transform 1 0 9844 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 1723858470
transform 1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1723858470
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_125
timestamp 1723858470
transform 1 0 12052 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_133
timestamp 1723858470
transform 1 0 12788 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_163
timestamp 1723858470
transform 1 0 15548 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1723858470
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_177
timestamp 1723858470
transform 1 0 16836 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_189
timestamp 1723858470
transform 1 0 17940 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_197
timestamp 1723858470
transform 1 0 18676 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_201
timestamp 1723858470
transform 1 0 19044 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_213
timestamp 1723858470
transform 1 0 20148 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 1723858470
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_225
timestamp 1723858470
transform 1 0 21252 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_232
timestamp 1723858470
transform 1 0 21896 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_244
timestamp 1723858470
transform 1 0 23000 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1723858470
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1723858470
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1723858470
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_29
timestamp 1723858470
transform 1 0 3220 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_37
timestamp 1723858470
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_63
timestamp 1723858470
transform 1 0 6348 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_85
timestamp 1723858470
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_113
timestamp 1723858470
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_131
timestamp 1723858470
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_146
timestamp 1723858470
transform 1 0 13984 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_154
timestamp 1723858470
transform 1 0 14720 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_185
timestamp 1723858470
transform 1 0 17572 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_189
timestamp 1723858470
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_213
timestamp 1723858470
transform 1 0 20148 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_225
timestamp 1723858470
transform 1 0 21252 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_233
timestamp 1723858470
transform 1 0 21988 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_242
timestamp 1723858470
transform 1 0 22816 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1723858470
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1723858470
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_27
timestamp 1723858470
transform 1 0 3036 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_47
timestamp 1723858470
transform 1 0 4876 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1723858470
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_70
timestamp 1723858470
transform 1 0 6992 0 -1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_77
timestamp 1723858470
transform 1 0 7636 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_89
timestamp 1723858470
transform 1 0 8740 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_96
timestamp 1723858470
transform 1 0 9384 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_104
timestamp 1723858470
transform 1 0 10120 0 -1 17952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1723858470
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1723858470
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1723858470
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1723858470
transform 1 0 14260 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1723858470
transform 1 0 15364 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1723858470
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_177
timestamp 1723858470
transform 1 0 16836 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_212
timestamp 1723858470
transform 1 0 20056 0 -1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1723858470
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1723858470
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1723858470
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_29
timestamp 1723858470
transform 1 0 3220 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_37
timestamp 1723858470
transform 1 0 3956 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_63
timestamp 1723858470
transform 1 0 6348 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_72
timestamp 1723858470
transform 1 0 7176 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1723858470
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_93
timestamp 1723858470
transform 1 0 9108 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_105
timestamp 1723858470
transform 1 0 10212 0 1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_126
timestamp 1723858470
transform 1 0 12144 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1723858470
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_141
timestamp 1723858470
transform 1 0 13524 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_157
timestamp 1723858470
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_164
timestamp 1723858470
transform 1 0 15640 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_176
timestamp 1723858470
transform 1 0 16744 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_182
timestamp 1723858470
transform 1 0 17296 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1723858470
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_211
timestamp 1723858470
transform 1 0 19964 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_223
timestamp 1723858470
transform 1 0 21068 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1723858470
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1723858470
transform 1 0 1932 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1723858470
transform 1 0 3036 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_39
timestamp 1723858470
transform 1 0 4140 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_47
timestamp 1723858470
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_54
timestamp 1723858470
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_57
timestamp 1723858470
transform 1 0 5796 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_81
timestamp 1723858470
transform 1 0 8004 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_104
timestamp 1723858470
transform 1 0 10120 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_133
timestamp 1723858470
transform 1 0 12788 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_140
timestamp 1723858470
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_173
timestamp 1723858470
transform 1 0 16468 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_181
timestamp 1723858470
transform 1 0 17204 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_192
timestamp 1723858470
transform 1 0 18216 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_204
timestamp 1723858470
transform 1 0 19320 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_210
timestamp 1723858470
transform 1 0 19872 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_216
timestamp 1723858470
transform 1 0 20424 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_225
timestamp 1723858470
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1723858470
transform 1 0 828 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1723858470
transform 1 0 1932 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1723858470
transform 1 0 3036 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_29
timestamp 1723858470
transform 1 0 3220 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_37
timestamp 1723858470
transform 1 0 3956 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_57
timestamp 1723858470
transform 1 0 5796 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_65
timestamp 1723858470
transform 1 0 6532 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_69
timestamp 1723858470
transform 1 0 6900 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_93
timestamp 1723858470
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_117
timestamp 1723858470
transform 1 0 11316 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_157
timestamp 1723858470
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_169
timestamp 1723858470
transform 1 0 16100 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_173
timestamp 1723858470
transform 1 0 16468 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_184
timestamp 1723858470
transform 1 0 17480 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1723858470
transform 1 0 18492 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_200
timestamp 1723858470
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_218
timestamp 1723858470
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_243
timestamp 1723858470
transform 1 0 22908 0 1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1723858470
transform 1 0 828 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1723858470
transform 1 0 1932 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_27
timestamp 1723858470
transform 1 0 3036 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_35
timestamp 1723858470
transform 1 0 3772 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1723858470
transform 1 0 5612 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_64
timestamp 1723858470
transform 1 0 6440 0 -1 20128
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_73
timestamp 1723858470
transform 1 0 7268 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_85
timestamp 1723858470
transform 1 0 8372 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_89
timestamp 1723858470
transform 1 0 8740 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_147
timestamp 1723858470
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_159
timestamp 1723858470
transform 1 0 15180 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1723858470
transform 1 0 15916 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_169
timestamp 1723858470
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_183
timestamp 1723858470
transform 1 0 17388 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_197
timestamp 1723858470
transform 1 0 18676 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1723858470
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1723858470
transform 1 0 828 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1723858470
transform 1 0 1932 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1723858470
transform 1 0 3036 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_29
timestamp 1723858470
transform 1 0 3220 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_37
timestamp 1723858470
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_50
timestamp 1723858470
transform 1 0 5152 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_61
timestamp 1723858470
transform 1 0 6164 0 1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_70
timestamp 1723858470
transform 1 0 6992 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_82
timestamp 1723858470
transform 1 0 8096 0 1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1723858470
transform 1 0 8372 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_97
timestamp 1723858470
transform 1 0 9476 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_103
timestamp 1723858470
transform 1 0 10028 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_111
timestamp 1723858470
transform 1 0 10764 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_119
timestamp 1723858470
transform 1 0 11500 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_127
timestamp 1723858470
transform 1 0 12236 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_135
timestamp 1723858470
transform 1 0 12972 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1723858470
transform 1 0 13340 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1723858470
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1723858470
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1723858470
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1723858470
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1723858470
transform 1 0 17940 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1723858470
transform 1 0 18492 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_197
timestamp 1723858470
transform 1 0 18676 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_207
timestamp 1723858470
transform 1 0 19596 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_215
timestamp 1723858470
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_240
timestamp 1723858470
transform 1 0 22632 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_244
timestamp 1723858470
transform 1 0 23000 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1723858470
transform 1 0 828 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1723858470
transform 1 0 1932 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1723858470
transform 1 0 3036 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1723858470
transform 1 0 4140 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_51
timestamp 1723858470
transform 1 0 5244 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_64
timestamp 1723858470
transform 1 0 6440 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_80
timestamp 1723858470
transform 1 0 7912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_100
timestamp 1723858470
transform 1 0 9752 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_109
timestamp 1723858470
transform 1 0 10580 0 -1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1723858470
transform 1 0 10948 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1723858470
transform 1 0 12052 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_137
timestamp 1723858470
transform 1 0 13156 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_153
timestamp 1723858470
transform 1 0 14628 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_161
timestamp 1723858470
transform 1 0 15364 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_172
timestamp 1723858470
transform 1 0 16376 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_176
timestamp 1723858470
transform 1 0 16744 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_184
timestamp 1723858470
transform 1 0 17480 0 -1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_191
timestamp 1723858470
transform 1 0 18124 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_203
timestamp 1723858470
transform 1 0 19228 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_211
timestamp 1723858470
transform 1 0 19964 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_232
timestamp 1723858470
transform 1 0 21896 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_244
timestamp 1723858470
transform 1 0 23000 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1723858470
transform 1 0 828 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1723858470
transform 1 0 1932 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1723858470
transform 1 0 3036 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_29
timestamp 1723858470
transform 1 0 3220 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_37
timestamp 1723858470
transform 1 0 3956 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_75
timestamp 1723858470
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_107
timestamp 1723858470
transform 1 0 10396 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_154
timestamp 1723858470
transform 1 0 14720 0 1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_200
timestamp 1723858470
transform 1 0 18952 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_231
timestamp 1723858470
transform 1 0 21804 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_243
timestamp 1723858470
transform 1 0 22908 0 1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1723858470
transform 1 0 828 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1723858470
transform 1 0 1932 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1723858470
transform 1 0 3036 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_39
timestamp 1723858470
transform 1 0 4140 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_43
timestamp 1723858470
transform 1 0 4508 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_54
timestamp 1723858470
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_153
timestamp 1723858470
transform 1 0 14628 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_191
timestamp 1723858470
transform 1 0 18124 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1723858470
transform 1 0 21068 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_241
timestamp 1723858470
transform 1 0 22724 0 -1 22304
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1723858470
transform 1 0 828 0 1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1723858470
transform 1 0 1932 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1723858470
transform 1 0 3036 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1723858470
transform 1 0 3220 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_41
timestamp 1723858470
transform 1 0 4324 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_85
timestamp 1723858470
transform 1 0 8372 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_107
timestamp 1723858470
transform 1 0 10396 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_117
timestamp 1723858470
transform 1 0 11316 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_125
timestamp 1723858470
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_138
timestamp 1723858470
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_151
timestamp 1723858470
transform 1 0 14444 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_159
timestamp 1723858470
transform 1 0 15180 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_165
timestamp 1723858470
transform 1 0 15732 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_210
timestamp 1723858470
transform 1 0 19872 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_236
timestamp 1723858470
transform 1 0 22264 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_244
timestamp 1723858470
transform 1 0 23000 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_3
timestamp 1723858470
transform 1 0 828 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_11
timestamp 1723858470
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_16
timestamp 1723858470
transform 1 0 2024 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_29
timestamp 1723858470
transform 1 0 3220 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_41
timestamp 1723858470
transform 1 0 4324 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_45
timestamp 1723858470
transform 1 0 4692 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1723858470
transform 1 0 5428 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_68
timestamp 1723858470
transform 1 0 6808 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_76
timestamp 1723858470
transform 1 0 7544 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_80
timestamp 1723858470
transform 1 0 7912 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_85
timestamp 1723858470
transform 1 0 8372 0 -1 23392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1723858470
transform 1 0 9108 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1723858470
transform 1 0 10212 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1723858470
transform 1 0 10764 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_119
timestamp 1723858470
transform 1 0 11500 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_131
timestamp 1723858470
transform 1 0 12604 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_139
timestamp 1723858470
transform 1 0 13340 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_147
timestamp 1723858470
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_159
timestamp 1723858470
transform 1 0 15180 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1723858470
transform 1 0 15916 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_169
timestamp 1723858470
transform 1 0 16100 0 -1 23392
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_176
timestamp 1723858470
transform 1 0 16744 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_188
timestamp 1723858470
transform 1 0 17848 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_211
timestamp 1723858470
transform 1 0 19964 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_217
timestamp 1723858470
transform 1 0 20516 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1723858470
transform 1 0 21068 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_230
timestamp 1723858470
transform 1 0 21712 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_236
timestamp 1723858470
transform 1 0 22264 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_243
timestamp 1723858470
transform 1 0 22908 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1723858470
transform -1 0 23092 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 22816 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1723858470
transform 1 0 1748 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1723858470
transform 1 0 5152 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1723858470
transform -1 0 7912 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1723858470
transform 1 0 10948 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 13524 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1723858470
transform 1 0 16468 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1723858470
transform 1 0 19412 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1723858470
transform 1 0 22356 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_42
timestamp 1723858470
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1723858470
transform -1 0 23368 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_43
timestamp 1723858470
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1723858470
transform -1 0 23368 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_44
timestamp 1723858470
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1723858470
transform -1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_45
timestamp 1723858470
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1723858470
transform -1 0 23368 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_46
timestamp 1723858470
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1723858470
transform -1 0 23368 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_47
timestamp 1723858470
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1723858470
transform -1 0 23368 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_48
timestamp 1723858470
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1723858470
transform -1 0 23368 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_49
timestamp 1723858470
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1723858470
transform -1 0 23368 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_50
timestamp 1723858470
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1723858470
transform -1 0 23368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_51
timestamp 1723858470
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1723858470
transform -1 0 23368 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_52
timestamp 1723858470
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1723858470
transform -1 0 23368 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_53
timestamp 1723858470
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1723858470
transform -1 0 23368 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_54
timestamp 1723858470
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1723858470
transform -1 0 23368 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_55
timestamp 1723858470
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1723858470
transform -1 0 23368 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_56
timestamp 1723858470
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1723858470
transform -1 0 23368 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_57
timestamp 1723858470
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1723858470
transform -1 0 23368 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_58
timestamp 1723858470
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1723858470
transform -1 0 23368 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_59
timestamp 1723858470
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1723858470
transform -1 0 23368 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_60
timestamp 1723858470
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1723858470
transform -1 0 23368 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_61
timestamp 1723858470
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1723858470
transform -1 0 23368 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_62
timestamp 1723858470
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1723858470
transform -1 0 23368 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_63
timestamp 1723858470
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1723858470
transform -1 0 23368 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_64
timestamp 1723858470
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1723858470
transform -1 0 23368 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_65
timestamp 1723858470
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1723858470
transform -1 0 23368 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_66
timestamp 1723858470
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1723858470
transform -1 0 23368 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_67
timestamp 1723858470
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1723858470
transform -1 0 23368 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_68
timestamp 1723858470
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1723858470
transform -1 0 23368 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_69
timestamp 1723858470
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1723858470
transform -1 0 23368 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_70
timestamp 1723858470
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1723858470
transform -1 0 23368 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_71
timestamp 1723858470
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1723858470
transform -1 0 23368 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_72
timestamp 1723858470
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1723858470
transform -1 0 23368 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_73
timestamp 1723858470
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1723858470
transform -1 0 23368 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_74
timestamp 1723858470
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1723858470
transform -1 0 23368 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_75
timestamp 1723858470
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1723858470
transform -1 0 23368 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_76
timestamp 1723858470
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1723858470
transform -1 0 23368 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_77
timestamp 1723858470
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1723858470
transform -1 0 23368 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_78
timestamp 1723858470
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1723858470
transform -1 0 23368 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_79
timestamp 1723858470
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1723858470
transform -1 0 23368 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_80
timestamp 1723858470
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1723858470
transform -1 0 23368 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_81
timestamp 1723858470
transform 1 0 552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1723858470
transform -1 0 23368 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_82
timestamp 1723858470
transform 1 0 552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1723858470
transform -1 0 23368 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_83
timestamp 1723858470
transform 1 0 552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1723858470
transform -1 0 23368 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1723858470
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1723858470
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1723858470
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1723858470
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_89
timestamp 1723858470
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_90
timestamp 1723858470
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_91
timestamp 1723858470
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1723858470
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1723858470
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_94
timestamp 1723858470
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_95
timestamp 1723858470
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1723858470
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1723858470
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1723858470
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1723858470
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1723858470
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1723858470
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1723858470
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1723858470
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_104
timestamp 1723858470
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1723858470
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1723858470
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1723858470
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_108
timestamp 1723858470
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_109
timestamp 1723858470
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_110
timestamp 1723858470
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1723858470
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_112
timestamp 1723858470
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_113
timestamp 1723858470
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_114
timestamp 1723858470
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_115
timestamp 1723858470
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1723858470
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_117
timestamp 1723858470
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_118
timestamp 1723858470
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_119
timestamp 1723858470
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1723858470
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1723858470
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1723858470
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_123
timestamp 1723858470
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1723858470
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1723858470
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1723858470
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1723858470
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1723858470
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1723858470
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1723858470
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1723858470
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp 1723858470
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp 1723858470
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1723858470
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1723858470
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_136
timestamp 1723858470
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_137
timestamp 1723858470
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_138
timestamp 1723858470
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1723858470
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_140
timestamp 1723858470
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_141
timestamp 1723858470
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_142
timestamp 1723858470
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_143
timestamp 1723858470
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_144
timestamp 1723858470
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_145
timestamp 1723858470
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_146
timestamp 1723858470
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_147
timestamp 1723858470
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_148
timestamp 1723858470
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_149
timestamp 1723858470
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_150
timestamp 1723858470
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_151
timestamp 1723858470
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_152
timestamp 1723858470
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_153
timestamp 1723858470
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_154
timestamp 1723858470
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_155
timestamp 1723858470
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp 1723858470
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_157
timestamp 1723858470
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_158
timestamp 1723858470
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_159
timestamp 1723858470
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp 1723858470
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp 1723858470
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_162
timestamp 1723858470
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_163
timestamp 1723858470
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp 1723858470
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp 1723858470
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_166
timestamp 1723858470
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_167
timestamp 1723858470
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp 1723858470
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp 1723858470
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_170
timestamp 1723858470
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_171
timestamp 1723858470
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp 1723858470
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp 1723858470
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_174
timestamp 1723858470
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_175
timestamp 1723858470
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_176
timestamp 1723858470
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp 1723858470
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_178
timestamp 1723858470
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_179
timestamp 1723858470
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_180
timestamp 1723858470
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_181
timestamp 1723858470
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_182
timestamp 1723858470
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_183
timestamp 1723858470
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_184
timestamp 1723858470
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_185
timestamp 1723858470
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_186
timestamp 1723858470
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_187
timestamp 1723858470
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_188
timestamp 1723858470
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_189
timestamp 1723858470
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_190
timestamp 1723858470
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_191
timestamp 1723858470
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_192
timestamp 1723858470
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_193
timestamp 1723858470
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_194
timestamp 1723858470
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_195
timestamp 1723858470
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_196
timestamp 1723858470
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_197
timestamp 1723858470
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_198
timestamp 1723858470
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_199
timestamp 1723858470
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_200
timestamp 1723858470
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_201
timestamp 1723858470
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_202
timestamp 1723858470
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_203
timestamp 1723858470
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_204
timestamp 1723858470
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_205
timestamp 1723858470
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_206
timestamp 1723858470
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_207
timestamp 1723858470
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_208
timestamp 1723858470
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_209
timestamp 1723858470
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_210
timestamp 1723858470
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_211
timestamp 1723858470
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_212
timestamp 1723858470
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_213
timestamp 1723858470
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_214
timestamp 1723858470
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_215
timestamp 1723858470
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_216
timestamp 1723858470
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_217
timestamp 1723858470
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_218
timestamp 1723858470
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_219
timestamp 1723858470
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_220
timestamp 1723858470
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_221
timestamp 1723858470
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_222
timestamp 1723858470
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_223
timestamp 1723858470
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_224
timestamp 1723858470
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_225
timestamp 1723858470
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_226
timestamp 1723858470
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_227
timestamp 1723858470
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_228
timestamp 1723858470
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_229
timestamp 1723858470
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_230
timestamp 1723858470
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_231
timestamp 1723858470
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_232
timestamp 1723858470
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_233
timestamp 1723858470
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_234
timestamp 1723858470
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_235
timestamp 1723858470
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_236
timestamp 1723858470
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_237
timestamp 1723858470
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_238
timestamp 1723858470
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_239
timestamp 1723858470
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_240
timestamp 1723858470
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_241
timestamp 1723858470
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_242
timestamp 1723858470
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_243
timestamp 1723858470
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_244
timestamp 1723858470
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_245
timestamp 1723858470
transform 1 0 10856 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_246
timestamp 1723858470
transform 1 0 16008 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_247
timestamp 1723858470
transform 1 0 21160 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_248
timestamp 1723858470
transform 1 0 3128 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_249
timestamp 1723858470
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_250
timestamp 1723858470
transform 1 0 13432 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_251
timestamp 1723858470
transform 1 0 18584 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_252
timestamp 1723858470
transform 1 0 3128 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_253
timestamp 1723858470
transform 1 0 5704 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_254
timestamp 1723858470
transform 1 0 8280 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_255
timestamp 1723858470
transform 1 0 10856 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_256
timestamp 1723858470
transform 1 0 13432 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_257
timestamp 1723858470
transform 1 0 16008 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_258
timestamp 1723858470
transform 1 0 18584 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_259
timestamp 1723858470
transform 1 0 21160 0 -1 23392
box -38 -48 130 592
<< labels >>
flabel metal4 s 4316 496 4636 23440 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3656 496 3976 23440 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 23600 3816 24000 3936 0 FreeSans 480 0 0 0 clk_in
port 2 nsew signal input
flabel metal3 s 23600 19592 24000 19712 0 FreeSans 480 0 0 0 clk_out
port 3 nsew signal output
flabel metal3 s 23600 11704 24000 11824 0 FreeSans 480 0 0 0 nrst
port 4 nsew signal input
flabel metal2 s 1674 23600 1730 24000 0 FreeSans 224 90 0 0 scale[0]
port 5 nsew signal input
flabel metal2 s 4618 23600 4674 24000 0 FreeSans 224 90 0 0 scale[1]
port 6 nsew signal input
flabel metal2 s 7562 23600 7618 24000 0 FreeSans 224 90 0 0 scale[2]
port 7 nsew signal input
flabel metal2 s 10506 23600 10562 24000 0 FreeSans 224 90 0 0 scale[3]
port 8 nsew signal input
flabel metal2 s 13450 23600 13506 24000 0 FreeSans 224 90 0 0 scale[4]
port 9 nsew signal input
flabel metal2 s 16394 23600 16450 24000 0 FreeSans 224 90 0 0 scale[5]
port 10 nsew signal input
flabel metal2 s 19338 23600 19394 24000 0 FreeSans 224 90 0 0 scale[6]
port 11 nsew signal input
flabel metal2 s 22282 23600 22338 24000 0 FreeSans 224 90 0 0 scale[7]
port 12 nsew signal input
rlabel metal1 11960 23392 11960 23392 0 VGND
rlabel metal1 11960 22848 11960 22848 0 VPWR
rlabel metal1 5392 13838 5392 13838 0 _0000_
rlabel metal1 4400 14518 4400 14518 0 _0001_
rlabel metal1 4733 12342 4733 12342 0 _0002_
rlabel metal1 5331 12750 5331 12750 0 _0003_
rlabel metal1 6389 12682 6389 12682 0 _0004_
rlabel via1 8689 11662 8689 11662 0 _0005_
rlabel metal2 8694 10982 8694 10982 0 _0006_
rlabel metal1 11316 10778 11316 10778 0 _0007_
rlabel via1 10989 11662 10989 11662 0 _0008_
rlabel metal1 12185 12342 12185 12342 0 _0009_
rlabel metal1 13744 12750 13744 12750 0 _0010_
rlabel metal1 13795 11254 13795 11254 0 _0011_
rlabel via1 14669 11662 14669 11662 0 _0012_
rlabel metal1 15885 13430 15885 13430 0 _0013_
rlabel via1 15957 14926 15957 14926 0 _0014_
rlabel metal1 16601 14518 16601 14518 0 _0015_
rlabel metal1 18706 17034 18706 17034 0 _0016_
rlabel metal1 19841 17782 19841 17782 0 _0017_
rlabel metal1 19499 19210 19499 19210 0 _0018_
rlabel metal1 21328 17782 21328 17782 0 _0019_
rlabel metal2 22310 19006 22310 19006 0 _0020_
rlabel via1 21109 19278 21109 19278 0 _0021_
rlabel metal1 3848 5814 3848 5814 0 _0022_
rlabel metal1 5294 6222 5294 6222 0 _0023_
rlabel metal1 4360 6834 4360 6834 0 _0024_
rlabel metal1 4360 7310 4360 7310 0 _0025_
rlabel metal1 3997 9078 3997 9078 0 _0026_
rlabel via1 4273 9486 4273 9486 0 _0027_
rlabel metal2 6118 8806 6118 8806 0 _0028_
rlabel metal1 6930 7242 6930 7242 0 _0029_
rlabel metal1 8560 6834 8560 6834 0 _0030_
rlabel metal1 8735 7242 8735 7242 0 _0031_
rlabel metal1 11168 6834 11168 6834 0 _0032_
rlabel metal2 10258 7106 10258 7106 0 _0033_
rlabel via1 12470 7310 12470 7310 0 _0034_
rlabel metal1 13738 7242 13738 7242 0 _0035_
rlabel via1 14678 7990 14678 7990 0 _0036_
rlabel metal2 15042 8194 15042 8194 0 _0037_
rlabel metal2 16974 8058 16974 8058 0 _0038_
rlabel metal2 16790 9282 16790 9282 0 _0039_
rlabel via1 18266 10574 18266 10574 0 _0040_
rlabel metal1 18982 12342 18982 12342 0 _0041_
rlabel metal1 17940 12614 17940 12614 0 _0042_
rlabel via1 19729 12750 19729 12750 0 _0043_
rlabel metal1 19780 10778 19780 10778 0 _0044_
rlabel metal2 20930 13396 20930 13396 0 _0045_
rlabel metal2 22034 11798 22034 11798 0 _0046_
rlabel metal1 21650 11594 21650 11594 0 _0047_
rlabel metal1 21558 9418 21558 9418 0 _0048_
rlabel metal2 21206 8636 21206 8636 0 _0049_
rlabel metal1 21620 7514 21620 7514 0 _0050_
rlabel metal1 20097 7990 20097 7990 0 _0051_
rlabel metal2 18814 8194 18814 8194 0 _0052_
rlabel via1 18809 9078 18809 9078 0 _0053_
rlabel via1 21937 18122 21937 18122 0 _0054_
rlabel metal2 23046 18156 23046 18156 0 _0055_
rlabel metal1 21252 18938 21252 18938 0 _0056_
rlabel metal1 5290 16694 5290 16694 0 _0057_
rlabel metal2 4738 17408 4738 17408 0 _0058_
rlabel metal1 6946 20570 6946 20570 0 _0059_
rlabel metal1 20194 21862 20194 21862 0 _0060_
rlabel metal1 5520 10778 5520 10778 0 _0061_
rlabel metal1 7176 9894 7176 9894 0 _0062_
rlabel metal2 8602 9690 8602 9690 0 _0063_
rlabel metal1 12742 10608 12742 10608 0 _0064_
rlabel metal1 12696 10098 12696 10098 0 _0065_
rlabel metal1 13294 10676 13294 10676 0 _0066_
rlabel metal2 14214 10234 14214 10234 0 _0067_
rlabel metal1 16790 13294 16790 13294 0 _0068_
rlabel metal1 17112 14042 17112 14042 0 _0069_
rlabel metal1 19182 16048 19182 16048 0 _0070_
rlabel metal1 20332 15946 20332 15946 0 _0071_
rlabel metal2 21666 16218 21666 16218 0 _0072_
rlabel metal1 21942 14416 21942 14416 0 _0073_
rlabel metal1 22241 9894 22241 9894 0 _0074_
rlabel metal1 4370 15674 4370 15674 0 _0075_
rlabel metal1 5060 14926 5060 14926 0 _0076_
rlabel metal2 5106 20196 5106 20196 0 _0077_
rlabel metal1 5014 19686 5014 19686 0 _0078_
rlabel metal2 5198 19686 5198 19686 0 _0079_
rlabel via2 4830 19261 4830 19261 0 _0080_
rlabel metal1 4416 17306 4416 17306 0 _0081_
rlabel metal1 8326 20910 8326 20910 0 _0082_
rlabel metal1 6348 13498 6348 13498 0 _0083_
rlabel metal2 8510 18462 8510 18462 0 _0084_
rlabel metal2 9614 19822 9614 19822 0 _0085_
rlabel metal1 8142 22746 8142 22746 0 _0086_
rlabel metal1 6624 20774 6624 20774 0 _0087_
rlabel metal1 9384 21862 9384 21862 0 _0088_
rlabel metal1 9430 21012 9430 21012 0 _0089_
rlabel metal1 7406 23018 7406 23018 0 _0090_
rlabel metal1 8556 21454 8556 21454 0 _0091_
rlabel metal2 8326 17612 8326 17612 0 _0092_
rlabel metal1 8418 22406 8418 22406 0 _0093_
rlabel metal1 9016 18802 9016 18802 0 _0094_
rlabel metal1 6907 21386 6907 21386 0 _0095_
rlabel metal1 6256 18802 6256 18802 0 _0096_
rlabel metal1 4094 18224 4094 18224 0 _0097_
rlabel metal2 6578 18564 6578 18564 0 _0098_
rlabel metal1 8188 19210 8188 19210 0 _0099_
rlabel metal2 7498 19108 7498 19108 0 _0100_
rlabel metal1 8970 17850 8970 17850 0 _0101_
rlabel metal1 8970 18666 8970 18666 0 _0102_
rlabel metal1 9062 17748 9062 17748 0 _0103_
rlabel metal1 8050 14382 8050 14382 0 _0104_
rlabel metal2 8970 13838 8970 13838 0 _0105_
rlabel metal2 8418 14042 8418 14042 0 _0106_
rlabel metal1 8694 13838 8694 13838 0 _0107_
rlabel metal1 8924 13974 8924 13974 0 _0108_
rlabel metal1 8510 12750 8510 12750 0 _0109_
rlabel metal1 8188 13158 8188 13158 0 _0110_
rlabel metal1 11592 19890 11592 19890 0 _0111_
rlabel metal1 9982 15572 9982 15572 0 _0112_
rlabel metal1 10718 19924 10718 19924 0 _0113_
rlabel metal1 10258 18666 10258 18666 0 _0114_
rlabel metal2 5934 18428 5934 18428 0 _0115_
rlabel metal2 7406 17408 7406 17408 0 _0116_
rlabel metal1 7314 17204 7314 17204 0 _0117_
rlabel metal2 8878 17306 8878 17306 0 _0118_
rlabel metal1 9154 17136 9154 17136 0 _0119_
rlabel metal2 9522 17510 9522 17510 0 _0120_
rlabel metal1 9844 14450 9844 14450 0 _0121_
rlabel metal1 9568 13838 9568 13838 0 _0122_
rlabel metal2 8786 13566 8786 13566 0 _0123_
rlabel metal2 9154 12954 9154 12954 0 _0124_
rlabel metal2 9338 12954 9338 12954 0 _0125_
rlabel metal1 8970 12818 8970 12818 0 _0126_
rlabel metal1 9062 10642 9062 10642 0 _0127_
rlabel metal1 9844 17646 9844 17646 0 _0128_
rlabel metal1 7820 19822 7820 19822 0 _0129_
rlabel metal2 4738 16014 4738 16014 0 _0130_
rlabel metal2 6026 15300 6026 15300 0 _0131_
rlabel metal2 5658 17476 5658 17476 0 _0132_
rlabel metal2 6118 15232 6118 15232 0 _0133_
rlabel metal1 6762 15130 6762 15130 0 _0134_
rlabel metal1 7084 15470 7084 15470 0 _0135_
rlabel metal1 8878 15470 8878 15470 0 _0136_
rlabel metal1 8740 15470 8740 15470 0 _0137_
rlabel metal1 10074 14586 10074 14586 0 _0138_
rlabel metal2 9706 15198 9706 15198 0 _0139_
rlabel metal2 10074 14892 10074 14892 0 _0140_
rlabel metal1 9246 13736 9246 13736 0 _0141_
rlabel metal1 10258 13736 10258 13736 0 _0142_
rlabel metal2 9982 13804 9982 13804 0 _0143_
rlabel metal2 9798 12716 9798 12716 0 _0144_
rlabel metal1 9384 12682 9384 12682 0 _0145_
rlabel metal2 10902 11390 10902 11390 0 _0146_
rlabel metal1 15778 18836 15778 18836 0 _0147_
rlabel metal2 4692 20366 4692 20366 0 _0148_
rlabel metal2 7682 20978 7682 20978 0 _0149_
rlabel metal2 5290 17680 5290 17680 0 _0150_
rlabel metal2 5382 16252 5382 16252 0 _0151_
rlabel metal1 6072 15878 6072 15878 0 _0152_
rlabel metal1 6164 16082 6164 16082 0 _0153_
rlabel via1 7038 14926 7038 14926 0 _0154_
rlabel metal1 6946 14960 6946 14960 0 _0155_
rlabel metal1 12098 14824 12098 14824 0 _0156_
rlabel metal1 10534 15028 10534 15028 0 _0157_
rlabel metal1 12581 15130 12581 15130 0 _0158_
rlabel metal2 10350 14654 10350 14654 0 _0159_
rlabel via2 11454 14212 11454 14212 0 _0160_
rlabel metal1 9936 13838 9936 13838 0 _0161_
rlabel metal2 12742 14076 12742 14076 0 _0162_
rlabel metal2 10396 13838 10396 13838 0 _0163_
rlabel metal1 10442 13872 10442 13872 0 _0164_
rlabel metal1 11132 13906 11132 13906 0 _0165_
rlabel metal1 12558 14042 12558 14042 0 _0166_
rlabel metal2 11178 13260 11178 13260 0 _0167_
rlabel metal1 11408 12410 11408 12410 0 _0168_
rlabel metal1 16100 20842 16100 20842 0 _0169_
rlabel metal1 15640 22678 15640 22678 0 _0170_
rlabel metal1 15732 21522 15732 21522 0 _0171_
rlabel metal1 11040 21454 11040 21454 0 _0172_
rlabel metal1 16698 21590 16698 21590 0 _0173_
rlabel metal1 15134 21420 15134 21420 0 _0174_
rlabel metal1 7958 21488 7958 21488 0 _0175_
rlabel metal1 8142 21114 8142 21114 0 _0176_
rlabel metal1 10396 22542 10396 22542 0 _0177_
rlabel metal1 8832 21386 8832 21386 0 _0178_
rlabel metal2 10902 21964 10902 21964 0 _0179_
rlabel metal1 11408 16014 11408 16014 0 _0180_
rlabel metal1 9062 16082 9062 16082 0 _0181_
rlabel metal1 12374 15946 12374 15946 0 _0182_
rlabel metal1 11684 16082 11684 16082 0 _0183_
rlabel metal1 12650 14892 12650 14892 0 _0184_
rlabel metal1 12650 14790 12650 14790 0 _0185_
rlabel metal2 13202 14620 13202 14620 0 _0186_
rlabel metal2 13754 14620 13754 14620 0 _0187_
rlabel metal1 13110 13396 13110 13396 0 _0188_
rlabel metal2 12466 13430 12466 13430 0 _0189_
rlabel metal1 14076 12410 14076 12410 0 _0190_
rlabel metal1 13662 21454 13662 21454 0 _0191_
rlabel metal1 18860 22678 18860 22678 0 _0192_
rlabel metal1 18814 22066 18814 22066 0 _0193_
rlabel metal2 19182 22780 19182 22780 0 _0194_
rlabel via1 19734 21947 19734 21947 0 _0195_
rlabel metal2 12190 21726 12190 21726 0 _0196_
rlabel metal1 12604 22066 12604 22066 0 _0197_
rlabel metal1 12696 21454 12696 21454 0 _0198_
rlabel metal2 12834 22202 12834 22202 0 _0199_
rlabel metal1 12627 22542 12627 22542 0 _0200_
rlabel metal1 12972 21318 12972 21318 0 _0201_
rlabel metal1 13248 21522 13248 21522 0 _0202_
rlabel metal2 14398 21964 14398 21964 0 _0203_
rlabel metal1 13340 16014 13340 16014 0 _0204_
rlabel metal2 13018 15742 13018 15742 0 _0205_
rlabel metal1 13570 16218 13570 16218 0 _0206_
rlabel metal1 13708 14926 13708 14926 0 _0207_
rlabel metal2 13846 14144 13846 14144 0 _0208_
rlabel metal1 13616 13294 13616 13294 0 _0209_
rlabel metal2 13386 18972 13386 18972 0 _0210_
rlabel metal1 14260 21998 14260 21998 0 _0211_
rlabel metal2 12650 20128 12650 20128 0 _0212_
rlabel metal2 10442 21284 10442 21284 0 _0213_
rlabel metal1 11086 21386 11086 21386 0 _0214_
rlabel metal1 9384 22066 9384 22066 0 _0215_
rlabel metal1 11040 22610 11040 22610 0 _0216_
rlabel metal1 10987 22066 10987 22066 0 _0217_
rlabel metal1 12972 22134 12972 22134 0 _0218_
rlabel metal1 13432 21998 13432 21998 0 _0219_
rlabel metal1 14260 22202 14260 22202 0 _0220_
rlabel metal2 13846 21488 13846 21488 0 _0221_
rlabel metal2 13570 17119 13570 17119 0 _0222_
rlabel metal1 13662 16660 13662 16660 0 _0223_
rlabel metal1 13938 16592 13938 16592 0 _0224_
rlabel metal2 13570 15402 13570 15402 0 _0225_
rlabel metal1 14076 13838 14076 13838 0 _0226_
rlabel metal1 14076 14042 14076 14042 0 _0227_
rlabel metal1 14214 13974 14214 13974 0 _0228_
rlabel metal2 7866 20026 7866 20026 0 _0229_
rlabel metal1 9384 19278 9384 19278 0 _0230_
rlabel metal1 11822 20468 11822 20468 0 _0231_
rlabel metal2 12006 20842 12006 20842 0 _0232_
rlabel metal2 12558 19788 12558 19788 0 _0233_
rlabel metal2 13110 19652 13110 19652 0 _0234_
rlabel metal2 13018 19822 13018 19822 0 _0235_
rlabel metal2 13570 19516 13570 19516 0 _0236_
rlabel metal1 13869 19890 13869 19890 0 _0237_
rlabel metal1 13800 18802 13800 18802 0 _0238_
rlabel metal2 14030 18462 14030 18462 0 _0239_
rlabel metal2 14306 15504 14306 15504 0 _0240_
rlabel metal1 14398 16660 14398 16660 0 _0241_
rlabel metal1 14490 18258 14490 18258 0 _0242_
rlabel metal1 14950 12410 14950 12410 0 _0243_
rlabel via1 10442 18190 10442 18190 0 _0244_
rlabel metal2 10350 18938 10350 18938 0 _0245_
rlabel metal1 11224 18190 11224 18190 0 _0246_
rlabel via1 12006 18734 12006 18734 0 _0247_
rlabel metal2 12834 19108 12834 19108 0 _0248_
rlabel metal1 14582 19482 14582 19482 0 _0249_
rlabel metal1 14030 18938 14030 18938 0 _0250_
rlabel metal2 14214 19210 14214 19210 0 _0251_
rlabel metal1 14628 18394 14628 18394 0 _0252_
rlabel metal1 14214 18700 14214 18700 0 _0253_
rlabel metal1 15456 13838 15456 13838 0 _0254_
rlabel metal1 5566 18292 5566 18292 0 _0255_
rlabel metal2 6026 17612 6026 17612 0 _0256_
rlabel metal1 6946 18224 6946 18224 0 _0257_
rlabel metal2 6302 16898 6302 16898 0 _0258_
rlabel metal2 10258 16796 10258 16796 0 _0259_
rlabel metal1 10166 17102 10166 17102 0 _0260_
rlabel metal1 10994 17034 10994 17034 0 _0261_
rlabel metal1 11224 17170 11224 17170 0 _0262_
rlabel metal1 12788 17102 12788 17102 0 _0263_
rlabel metal2 12926 17646 12926 17646 0 _0264_
rlabel metal1 16606 17748 16606 17748 0 _0265_
rlabel metal2 16790 17306 16790 17306 0 _0266_
rlabel metal1 15594 16558 15594 16558 0 _0267_
rlabel metal2 15042 17884 15042 17884 0 _0268_
rlabel metal1 14950 16150 14950 16150 0 _0269_
rlabel metal1 15226 16558 15226 16558 0 _0270_
rlabel metal2 16330 15980 16330 15980 0 _0271_
rlabel metal2 16698 15708 16698 15708 0 _0272_
rlabel metal2 14950 21165 14950 21165 0 _0273_
rlabel metal1 5888 20366 5888 20366 0 _0274_
rlabel metal2 6026 20060 6026 20060 0 _0275_
rlabel metal2 6118 18938 6118 18938 0 _0276_
rlabel metal1 6762 19278 6762 19278 0 _0277_
rlabel metal1 6624 19754 6624 19754 0 _0278_
rlabel metal1 14766 18802 14766 18802 0 _0279_
rlabel metal1 14582 18734 14582 18734 0 _0280_
rlabel metal1 16008 18394 16008 18394 0 _0281_
rlabel metal1 15870 18768 15870 18768 0 _0282_
rlabel metal2 16514 18156 16514 18156 0 _0283_
rlabel metal1 14398 17170 14398 17170 0 _0284_
rlabel metal2 16330 17306 16330 17306 0 _0285_
rlabel metal1 16606 17170 16606 17170 0 _0286_
rlabel metal1 16008 16626 16008 16626 0 _0287_
rlabel metal1 16530 16694 16530 16694 0 _0288_
rlabel metal2 16974 15844 16974 15844 0 _0289_
rlabel metal1 17066 15572 17066 15572 0 _0290_
rlabel metal1 16146 21012 16146 21012 0 _0291_
rlabel metal1 17020 21658 17020 21658 0 _0292_
rlabel metal1 16560 20978 16560 20978 0 _0293_
rlabel metal1 17204 21454 17204 21454 0 _0294_
rlabel metal2 16698 21284 16698 21284 0 _0295_
rlabel metal1 16652 19890 16652 19890 0 _0296_
rlabel metal1 15088 19822 15088 19822 0 _0297_
rlabel metal1 17480 19958 17480 19958 0 _0298_
rlabel metal2 16882 19550 16882 19550 0 _0299_
rlabel metal1 17848 19686 17848 19686 0 _0300_
rlabel metal1 17802 18836 17802 18836 0 _0301_
rlabel metal1 17710 18768 17710 18768 0 _0302_
rlabel metal1 18492 18938 18492 18938 0 _0303_
rlabel metal2 17618 18394 17618 18394 0 _0304_
rlabel metal1 18446 18292 18446 18292 0 _0305_
rlabel metal1 14076 14586 14076 14586 0 _0306_
rlabel metal1 15272 16490 15272 16490 0 _0307_
rlabel metal1 17250 17034 17250 17034 0 _0308_
rlabel metal2 17158 17034 17158 17034 0 _0309_
rlabel metal1 17158 17136 17158 17136 0 _0310_
rlabel metal1 18308 17714 18308 17714 0 _0311_
rlabel metal1 18538 18394 18538 18394 0 _0312_
rlabel metal2 18354 17408 18354 17408 0 _0313_
rlabel metal1 18722 16762 18722 16762 0 _0314_
rlabel metal1 17664 21862 17664 21862 0 _0315_
rlabel metal1 17710 20978 17710 20978 0 _0316_
rlabel metal1 17802 21046 17802 21046 0 _0317_
rlabel metal1 18216 21522 18216 21522 0 _0318_
rlabel metal1 18538 21488 18538 21488 0 _0319_
rlabel via1 17810 19958 17810 19958 0 _0320_
rlabel metal2 18262 19482 18262 19482 0 _0321_
rlabel metal1 18400 19278 18400 19278 0 _0322_
rlabel metal2 17986 18700 17986 18700 0 _0323_
rlabel metal1 18768 18122 18768 18122 0 _0324_
rlabel metal1 19320 18190 19320 18190 0 _0325_
rlabel metal1 20792 22678 20792 22678 0 _0326_
rlabel metal2 21482 22950 21482 22950 0 _0327_
rlabel metal2 21206 22372 21206 22372 0 _0328_
rlabel metal1 21574 21930 21574 21930 0 _0329_
rlabel metal1 22218 22440 22218 22440 0 _0330_
rlabel metal2 21022 21658 21022 21658 0 _0331_
rlabel metal1 20470 21420 20470 21420 0 _0332_
rlabel metal1 20562 21522 20562 21522 0 _0333_
rlabel metal1 21252 21046 21252 21046 0 _0334_
rlabel metal2 20102 21148 20102 21148 0 _0335_
rlabel metal2 19550 20570 19550 20570 0 _0336_
rlabel metal1 18814 19958 18814 19958 0 _0337_
rlabel metal2 18722 19618 18722 19618 0 _0338_
rlabel metal2 18998 20094 18998 20094 0 _0339_
rlabel metal1 19642 19822 19642 19822 0 _0340_
rlabel metal2 19734 20060 19734 20060 0 _0341_
rlabel metal2 20010 19380 20010 19380 0 _0342_
rlabel metal2 21482 20196 21482 20196 0 _0343_
rlabel metal1 20838 21998 20838 21998 0 _0344_
rlabel metal2 22310 21760 22310 21760 0 _0345_
rlabel metal1 21528 21590 21528 21590 0 _0346_
rlabel metal1 21106 21114 21106 21114 0 _0347_
rlabel metal2 20654 20672 20654 20672 0 _0348_
rlabel metal1 20562 20400 20562 20400 0 _0349_
rlabel metal2 20930 18972 20930 18972 0 _0350_
rlabel metal1 21160 20434 21160 20434 0 _0351_
rlabel metal2 22678 19822 22678 19822 0 _0352_
rlabel metal1 21250 19890 21250 19890 0 _0353_
rlabel metal2 22770 9503 22770 9503 0 _0354_
rlabel metal1 22310 10234 22310 10234 0 _0355_
rlabel metal2 21850 15572 21850 15572 0 _0356_
rlabel metal1 22862 14484 22862 14484 0 _0357_
rlabel metal1 21298 9146 21298 9146 0 _0358_
rlabel metal2 22126 10336 22126 10336 0 _0359_
rlabel metal1 22678 14348 22678 14348 0 _0360_
rlabel metal1 22218 14926 22218 14926 0 _0361_
rlabel metal2 21482 15538 21482 15538 0 _0362_
rlabel metal1 21896 15062 21896 15062 0 _0363_
rlabel metal2 20746 15708 20746 15708 0 _0364_
rlabel metal2 20562 15130 20562 15130 0 _0365_
rlabel metal1 20792 15130 20792 15130 0 _0366_
rlabel metal2 19734 15708 19734 15708 0 _0367_
rlabel metal2 19734 15164 19734 15164 0 _0368_
rlabel metal1 20194 14994 20194 14994 0 _0369_
rlabel metal2 18630 14688 18630 14688 0 _0370_
rlabel metal1 19274 14382 19274 14382 0 _0371_
rlabel metal1 17902 14586 17902 14586 0 _0372_
rlabel metal1 18584 13838 18584 13838 0 _0373_
rlabel metal2 18722 14450 18722 14450 0 _0374_
rlabel metal2 19090 14144 19090 14144 0 _0375_
rlabel metal1 17304 13702 17304 13702 0 _0376_
rlabel metal1 18032 13430 18032 13430 0 _0377_
rlabel metal1 17848 13362 17848 13362 0 _0378_
rlabel metal1 18492 13498 18492 13498 0 _0379_
rlabel metal2 16698 11594 16698 11594 0 _0380_
rlabel metal2 16882 10778 16882 10778 0 _0381_
rlabel metal2 16238 10914 16238 10914 0 _0382_
rlabel metal1 16974 10778 16974 10778 0 _0383_
rlabel metal1 16698 10676 16698 10676 0 _0384_
rlabel metal2 14950 9758 14950 9758 0 _0385_
rlabel metal1 15594 9486 15594 9486 0 _0386_
rlabel metal2 14766 10268 14766 10268 0 _0387_
rlabel metal2 14490 9724 14490 9724 0 _0388_
rlabel metal1 15088 9690 15088 9690 0 _0389_
rlabel metal2 12466 10574 12466 10574 0 _0390_
rlabel metal2 13662 9996 13662 9996 0 _0391_
rlabel metal1 14858 9622 14858 9622 0 _0392_
rlabel metal2 11730 9418 11730 9418 0 _0393_
rlabel metal1 12558 8942 12558 8942 0 _0394_
rlabel metal1 12328 10098 12328 10098 0 _0395_
rlabel metal1 11914 9554 11914 9554 0 _0396_
rlabel metal2 12282 9078 12282 9078 0 _0397_
rlabel metal2 11086 9146 11086 9146 0 _0398_
rlabel metal1 11730 8874 11730 8874 0 _0399_
rlabel metal1 8862 10166 8862 10166 0 _0400_
rlabel metal1 9200 9010 9200 9010 0 _0401_
rlabel metal2 8234 9214 8234 9214 0 _0402_
rlabel metal2 8326 9248 8326 9248 0 _0403_
rlabel metal1 8786 8908 8786 8908 0 _0404_
rlabel via1 7322 10234 7322 10234 0 _0405_
rlabel metal2 7498 9690 7498 9690 0 _0406_
rlabel metal1 7682 9690 7682 9690 0 _0407_
rlabel metal1 5490 10506 5490 10506 0 _0408_
rlabel metal1 6578 10608 6578 10608 0 _0409_
rlabel metal1 6854 10778 6854 10778 0 _0410_
rlabel metal1 5566 11050 5566 11050 0 _0411_
rlabel metal2 6394 10404 6394 10404 0 _0412_
rlabel metal1 4738 7956 4738 7956 0 _0413_
rlabel metal2 3450 6800 3450 6800 0 _0414_
rlabel metal2 5474 7888 5474 7888 0 _0415_
rlabel metal1 5980 9690 5980 9690 0 _0416_
rlabel metal1 6056 9418 6056 9418 0 _0417_
rlabel metal1 5934 9588 5934 9588 0 _0418_
rlabel metal1 7268 9486 7268 9486 0 _0419_
rlabel metal1 8326 9078 8326 9078 0 _0420_
rlabel metal1 12282 9112 12282 9112 0 _0421_
rlabel metal1 14122 9146 14122 9146 0 _0422_
rlabel metal1 16284 9622 16284 9622 0 _0423_
rlabel metal1 18032 10438 18032 10438 0 _0424_
rlabel metal2 19458 14722 19458 14722 0 _0425_
rlabel metal1 21758 14926 21758 14926 0 _0426_
rlabel metal1 22126 14994 22126 14994 0 _0427_
rlabel metal2 22402 14518 22402 14518 0 _0428_
rlabel metal2 22034 18207 22034 18207 0 _0429_
rlabel metal1 21942 12818 21942 12818 0 _0430_
rlabel metal2 5658 7752 5658 7752 0 _0431_
rlabel metal1 3956 6426 3956 6426 0 _0432_
rlabel metal1 4232 6970 4232 6970 0 _0433_
rlabel metal2 3358 9792 3358 9792 0 _0434_
rlabel metal1 3726 9690 3726 9690 0 _0435_
rlabel metal2 6394 9792 6394 9792 0 _0436_
rlabel metal1 4600 9894 4600 9894 0 _0437_
rlabel metal1 5612 8534 5612 8534 0 _0438_
rlabel metal1 6072 8534 6072 8534 0 _0439_
rlabel metal2 6578 7616 6578 7616 0 _0440_
rlabel metal1 6808 6970 6808 6970 0 _0441_
rlabel metal1 7912 8058 7912 8058 0 _0442_
rlabel metal2 7866 7990 7866 7990 0 _0443_
rlabel metal1 9016 7786 9016 7786 0 _0444_
rlabel metal1 8924 7718 8924 7718 0 _0445_
rlabel metal1 10074 7752 10074 7752 0 _0446_
rlabel metal1 10396 6426 10396 6426 0 _0447_
rlabel metal2 10902 7684 10902 7684 0 _0448_
rlabel metal2 10442 7174 10442 7174 0 _0449_
rlabel via1 14590 8330 14590 8330 0 _0450_
rlabel metal1 12052 7718 12052 7718 0 _0451_
rlabel metal2 13202 7888 13202 7888 0 _0452_
rlabel metal1 13294 6970 13294 6970 0 _0453_
rlabel metal2 14766 7786 14766 7786 0 _0454_
rlabel metal1 13708 8058 13708 8058 0 _0455_
rlabel metal1 18078 8432 18078 8432 0 _0456_
rlabel metal2 15410 7616 15410 7616 0 _0457_
rlabel metal1 17572 7718 17572 7718 0 _0458_
rlabel metal1 17004 7990 17004 7990 0 _0459_
rlabel metal1 17664 8874 17664 8874 0 _0460_
rlabel metal1 16974 8840 16974 8840 0 _0461_
rlabel via1 18454 13430 18454 13430 0 _0462_
rlabel metal1 18078 10234 18078 10234 0 _0463_
rlabel metal1 17250 12070 17250 12070 0 _0464_
rlabel metal1 17848 11866 17848 11866 0 _0465_
rlabel metal1 19274 13226 19274 13226 0 _0466_
rlabel metal1 18400 12954 18400 12954 0 _0467_
rlabel metal1 20608 13226 20608 13226 0 _0468_
rlabel metal1 19780 11866 19780 11866 0 _0469_
rlabel metal1 20378 10778 20378 10778 0 _0470_
rlabel via1 20002 10506 20002 10506 0 _0471_
rlabel metal1 22205 11322 22205 11322 0 _0472_
rlabel metal2 21114 13056 21114 13056 0 _0473_
rlabel metal1 21620 11186 21620 11186 0 _0474_
rlabel metal1 21896 10982 21896 10982 0 _0475_
rlabel metal1 21328 10506 21328 10506 0 _0476_
rlabel metal2 21298 12546 21298 12546 0 _0477_
rlabel metal2 20746 9894 20746 9894 0 _0478_
rlabel metal1 21298 9690 21298 9690 0 _0479_
rlabel metal1 21344 8262 21344 8262 0 _0480_
rlabel metal1 22310 8330 22310 8330 0 _0481_
rlabel metal1 21160 7310 21160 7310 0 _0482_
rlabel metal1 21114 8330 21114 8330 0 _0483_
rlabel metal1 18630 8330 18630 8330 0 _0484_
rlabel metal1 18584 7990 18584 7990 0 _0485_
rlabel metal1 19504 7922 19504 7922 0 _0486_
rlabel metal1 19136 9690 19136 9690 0 _0487_
rlabel metal2 19550 8704 19550 8704 0 _0488_
rlabel metal1 21850 18156 21850 18156 0 _0489_
rlabel metal2 22954 3927 22954 3927 0 clk_in
rlabel metal2 23046 19737 23046 19737 0 clk_out
rlabel metal2 5842 7038 5842 7038 0 count\[0\]
rlabel metal1 11822 8330 11822 8330 0 count\[10\]
rlabel metal1 11224 8602 11224 8602 0 count\[11\]
rlabel metal1 11730 8398 11730 8398 0 count\[12\]
rlabel metal1 14444 8330 14444 8330 0 count\[13\]
rlabel metal1 13432 7786 13432 7786 0 count\[14\]
rlabel metal1 15088 8534 15088 8534 0 count\[15\]
rlabel metal2 17802 10676 17802 10676 0 count\[16\]
rlabel metal2 16698 10166 16698 10166 0 count\[17\]
rlabel metal1 17986 13872 17986 13872 0 count\[18\]
rlabel metal1 19136 12614 19136 12614 0 count\[19\]
rlabel metal2 6026 7038 6026 7038 0 count\[1\]
rlabel metal1 18492 13158 18492 13158 0 count\[20\]
rlabel metal2 20470 14110 20470 14110 0 count\[21\]
rlabel metal1 21022 15504 21022 15504 0 count\[22\]
rlabel metal1 21574 12954 21574 12954 0 count\[23\]
rlabel metal1 21712 13362 21712 13362 0 count\[24\]
rlabel metal1 22632 11526 22632 11526 0 count\[25\]
rlabel metal1 22402 10030 22402 10030 0 count\[26\]
rlabel metal2 22586 10336 22586 10336 0 count\[27\]
rlabel metal1 22724 8330 22724 8330 0 count\[28\]
rlabel metal1 22586 8534 22586 8534 0 count\[29\]
rlabel metal1 5934 6970 5934 6970 0 count\[2\]
rlabel metal1 20562 8942 20562 8942 0 count\[30\]
rlabel metal1 19591 9486 19591 9486 0 count\[31\]
rlabel via1 5566 6902 5566 6902 0 count\[3\]
rlabel metal1 6210 9486 6210 9486 0 count\[4\]
rlabel metal1 5198 9690 5198 9690 0 count\[5\]
rlabel metal1 5244 9078 5244 9078 0 count\[6\]
rlabel metal1 7866 10064 7866 10064 0 count\[7\]
rlabel metal2 7958 8704 7958 8704 0 count\[8\]
rlabel metal1 8418 7888 8418 7888 0 count\[9\]
rlabel metal2 22770 5712 22770 5712 0 net1
rlabel metal2 22678 22610 22678 22610 0 net10
rlabel metal1 7866 7956 7866 7956 0 net11
rlabel metal1 19826 13362 19826 13362 0 net12
rlabel metal1 13708 8262 13708 8262 0 net13
rlabel metal2 20746 8653 20746 8653 0 net14
rlabel metal1 14168 13362 14168 13362 0 net15
rlabel metal2 15226 14484 15226 14484 0 net16
rlabel metal1 15134 20978 15134 20978 0 net17
rlabel metal1 4784 19958 4784 19958 0 net18
rlabel metal1 4692 15538 4692 15538 0 net19
rlabel metal2 22862 11599 22862 11599 0 net2
rlabel metal1 5428 14926 5428 14926 0 net20
rlabel metal1 16284 15538 16284 15538 0 net21
rlabel metal2 20930 16150 20930 16150 0 net22
rlabel metal1 8694 7310 8694 7310 0 net23
rlabel metal1 4554 12716 4554 12716 0 net24
rlabel metal1 12742 7276 12742 7276 0 net25
rlabel metal1 23414 12036 23414 12036 0 net26
rlabel metal2 13570 12585 13570 12585 0 net27
rlabel metal1 16054 14382 16054 14382 0 net28
rlabel metal1 20378 13974 20378 13974 0 net29
rlabel metal1 1978 23086 1978 23086 0 net3
rlabel metal1 4370 20366 4370 20366 0 net4
rlabel metal2 5658 20672 5658 20672 0 net5
rlabel metal2 18170 22780 18170 22780 0 net6
rlabel metal2 20286 22882 20286 22882 0 net7
rlabel metal1 16974 22440 16974 22440 0 net8
rlabel metal2 22126 22304 22126 22304 0 net9
rlabel metal2 23046 11169 23046 11169 0 nrst
rlabel metal2 1794 23443 1794 23443 0 scale[0]
rlabel metal1 5198 23188 5198 23188 0 scale[1]
rlabel metal2 7866 23443 7866 23443 0 scale[2]
rlabel metal1 10810 23222 10810 23222 0 scale[3]
rlabel metal2 13570 23443 13570 23443 0 scale[4]
rlabel metal2 16514 23443 16514 23443 0 scale[5]
rlabel metal2 19412 23154 19412 23154 0 scale[6]
rlabel metal1 22356 23154 22356 23154 0 scale[7]
rlabel metal1 22724 18802 22724 18802 0 signal_clk_out
rlabel metal1 9200 11866 9200 11866 0 true_scale\[10\]
rlabel metal1 9568 10642 9568 10642 0 true_scale\[11\]
rlabel metal1 12926 10540 12926 10540 0 true_scale\[12\]
rlabel metal1 11914 11866 11914 11866 0 true_scale\[13\]
rlabel metal2 12006 12580 12006 12580 0 true_scale\[14\]
rlabel metal1 14720 12274 14720 12274 0 true_scale\[15\]
rlabel metal1 14582 11322 14582 11322 0 true_scale\[16\]
rlabel metal1 15456 11866 15456 11866 0 true_scale\[17\]
rlabel metal1 15594 13770 15594 13770 0 true_scale\[18\]
rlabel metal1 16974 15130 16974 15130 0 true_scale\[19\]
rlabel metal1 17526 14926 17526 14926 0 true_scale\[20\]
rlabel metal2 19274 16490 19274 16490 0 true_scale\[21\]
rlabel metal2 18630 17952 18630 17952 0 true_scale\[22\]
rlabel metal2 20378 18972 20378 18972 0 true_scale\[23\]
rlabel metal1 21298 17544 21298 17544 0 true_scale\[24\]
rlabel metal1 22678 18938 22678 18938 0 true_scale\[25\]
rlabel metal2 22218 19584 22218 19584 0 true_scale\[26\]
rlabel metal1 6118 13974 6118 13974 0 true_scale\[5\]
rlabel metal1 4738 14824 4738 14824 0 true_scale\[6\]
rlabel metal1 5474 12410 5474 12410 0 true_scale\[7\]
rlabel metal1 6072 12954 6072 12954 0 true_scale\[8\]
rlabel metal1 7130 12342 7130 12342 0 true_scale\[9\]
flabel metal4 3760 23520 3860 23600 0 FreeSans 320 0 0 0 VPWR
flabel metal4 4420 360 4520 420 0 FreeSans 320 0 0 0 VGND
<< properties >>
string FIXED_BBOX 0 0 24000 24000
<< end >>
