* NGSPICE file created from tt_um_hugodiasg_temp_sensor_clock_divider.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_FRXWNM a_n100_n297# a_100_n200# w_n194_n300# a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n194_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_FVXEPM a_n100_n297# a_100_n200# w_n194_n300# a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n194_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_FVTXNM a_29_n297# a_n287_n200# a_n229_n297# a_229_n200#
+ a_n29_n200# w_n323_n300#
X0 a_229_n200# a_29_n297# a_n29_n200# w_n323_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X1 a_n29_n200# a_n229_n297# a_n287_n200# w_n323_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_3HGYVM a_n100_n297# a_100_n200# w_n194_n300# a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n194_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_SKTYVM a_n500_n297# a_500_n200# w_n594_n300# a_n558_n200#
X0 a_500_n200# a_n500_n297# a_n558_n200# w_n594_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=5
.ends

.subckt sky130_fd_pr__nfet_01v8_9VJR3B a_100_527# a_n158_n727# a_100_n309# a_n100_21#
+ a_n158_n309# a_100_109# a_n158_527# a_n100_n815# a_n100_439# a_n158_109# a_100_n727#
+ a_n100_n397# VSUBS
X0 a_100_n309# a_n100_n397# a_n158_n309# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_527# a_n100_439# a_n158_527# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_n727# a_n100_n815# a_n158_n727# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_109# a_n100_21# a_n158_109# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_YAWWFM a_29_n297# a_n287_n200# w_n581_n300# a_n229_n297#
+ a_287_n297# a_229_n200# a_n545_n200# a_n487_n297# a_487_n200# a_n29_n200#
X0 a_229_n200# a_29_n297# a_n29_n200# w_n581_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_n29_n200# a_n229_n297# a_n287_n200# w_n581_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_n287_n200# a_n487_n297# a_n545_n200# w_n581_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X3 a_487_n200# a_287_n297# a_229_n200# w_n581_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_YAEUFM a_29_n297# a_n287_n200# a_n1061_n200# a_n745_n297#
+ a_745_n200# a_803_n297# a_n229_n297# a_n1003_n297# a_287_n297# a_229_n200# a_n545_n200#
+ a_1003_n200# a_n487_n297# a_487_n200# a_n29_n200# a_545_n297# a_n803_n200# w_n1097_n300#
X0 a_229_n200# a_29_n297# a_n29_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_n29_n200# a_n229_n297# a_n287_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_n545_n200# a_n745_n297# a_n803_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_n287_n200# a_n487_n297# a_n545_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_n803_n200# a_n1003_n297# a_n1061_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X5 a_1003_n200# a_803_n297# a_745_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X6 a_745_n200# a_545_n297# a_487_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_487_n200# a_287_n297# a_229_n200# w_n1097_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sensor vd vts vtd gnd
Xsky130_fd_pr__pfet_01v8_FRXWNM_0 vd vd vd vd sky130_fd_pr__pfet_01v8_FRXWNM
Xsky130_fd_pr__pfet_01v8_FRXWNM_1 vd vd vd vd sky130_fd_pr__pfet_01v8_FRXWNM
Xsky130_fd_pr__pfet_01v8_FRXWNM_2 vd vd vd vd sky130_fd_pr__pfet_01v8_FRXWNM
Xsky130_fd_pr__pfet_01v8_FRXWNM_3 vts vts vts vts sky130_fd_pr__pfet_01v8_FRXWNM
Xsky130_fd_pr__pfet_01v8_FVXEPM_0 c c vd c sky130_fd_pr__pfet_01v8_FVXEPM
Xsky130_fd_pr__pfet_01v8_FRXWNM_4 vts vts vts vts sky130_fd_pr__pfet_01v8_FRXWNM
XXP1 a a a a vd vd sky130_fd_pr__pfet_01v8_FVTXNM
XXP3 vtd d vd vd sky130_fd_pr__pfet_01v8_3HGYVM
XXP4 vtd vd vd vts sky130_fd_pr__pfet_01v8_SKTYVM
Xsky130_fd_pr__nfet_01v8_9VJR3B_0 gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd
+ gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_1 gnd a gnd b a gnd a b b a gnd b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_2 a gnd a b gnd a gnd b b gnd a b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_3 gnd vtd gnd b vtd gnd vtd b b vtd gnd b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_4 vtd gnd vtd b gnd vtd gnd b b gnd vtd b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_5 gnd b gnd b b gnd b b b b gnd b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_6 gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd
+ gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__nfet_01v8_9VJR3B_7 b gnd b b gnd b gnd b b gnd b b gnd sky130_fd_pr__nfet_01v8_9VJR3B
Xsky130_fd_pr__pfet_01v8_YAWWFM_0 a d vd a a d c a c c sky130_fd_pr__pfet_01v8_YAWWFM
Xsky130_fd_pr__pfet_01v8_YAWWFM_1 vtd b vd vtd vtd b c vtd c c sky130_fd_pr__pfet_01v8_YAWWFM
Xsky130_fd_pr__pfet_01v8_YAEUFM_0 vtd vts vtd vtd vts vtd vtd vtd vtd vts vtd vtd
+ vtd vtd vtd vtd vts vts sky130_fd_pr__pfet_01v8_YAEUFM
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X18 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 VPB VNB VGND VPWR A Y B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VPB VNB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB B C A X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_1 VPB VNB VGND VPWR A_N B Y
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VPB VNB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_4 VPB VNB VPWR VGND B C A X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.26 ps=1.45 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.20475 pd=1.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X5 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_109_297# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR VPB VNB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__a21boi_2 VNB VPB VPWR VGND B1_N A2 Y A1
X0 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183125 ps=1.24 w=0.65 l=0.15
X1 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_479_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 Y a_61_47# a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_61_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VGND A2 a_637_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_61_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A1 a_479_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.06825 ps=0.86 w=0.65 l=0.15
X11 VGND B1_N a_61_47# VNB sky130_fd_pr__nfet_01v8 ad=0.183125 pd=1.24 as=0.126 ps=1.44 w=0.42 l=0.15
X12 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X13 a_637_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 VPWR VGND VPB VNB B1_N Y A1 A2
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 VNB VPB VPWR VGND A X B
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 VPB VNB VGND VPWR X A B
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.91 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_2 VPWR VGND X B A VPB VNB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 B1 Y A1 VPB VNB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 VPB VNB VGND VPWR A B Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VPB VNB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VPB VNB
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.099125 ps=0.955 w=0.65 l=0.15
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 B2
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 VPB VNB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND VPB VNB A2 A1 B1 X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_1 VPB VNB VGND VPWR A1 Y C1 B1 A2
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.17225 ps=1.83 w=0.65 l=0.15
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0.39325 pd=2.51 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 VPB VNB X A3 A2 A1 B1 VGND VPWR
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 VPWR VGND VPB VNB B C A X D_N
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_1 VPWR VGND VPB VNB Y C1 B1 A1 A2
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 X A1 A2 A3 B1 VPB VNB VGND VPWR
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 X C A B D VGND VPWR VPB VNB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_2 VNB VPB VPWR VGND B1 Y A1 A2 A3
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X4 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
X11 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X13 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X14 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_2 VNB VPB VGND VPWR A2 A1 Y B1
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_2 VGND VPWR B1 A1 Y A2 VPB VNB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_4 VNB VPB VPWR VGND B1 Y A1 A2
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_2 VNB VPB VGND VPWR Y B1 A2 A1 C1
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_1 VNB VPB VGND VPWR X A2 A1 B1_N
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258375 ps=1.445 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258375 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 VGND VPWR VPB VNB B C A X
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB X A1 S A0
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 VNB VPB VGND VPWR X A2 B1 A1 C1
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 VNB VPB VGND VPWR B1_N A1 A2 X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_1 VPB VNB VPWR VGND A1 B1_N Y A2
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1275 pd=1.255 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1275 ps=1.255 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17825 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.17825 ps=1.4 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_4 VNB VPB VGND VPWR Y B A
X0 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X36 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_4 VNB VPB VGND VPWR B X A
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27245 ps=2.56 w=1 l=0.15
X15 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17875 ps=1.85 w=0.65 l=0.15
X17 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X19 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X24 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2568 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X30 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X38 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 VPB VNB VGND VPWR A B Y C
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 VNB VPB VGND VPWR X A1 A2 B1 C1
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_2 VNB VPB VGND VPWR A2 A1 B1 X
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1105 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1625 pd=1.15 as=0.1105 ps=0.99 w=0.65 l=0.15
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.1625 ps=1.15 w=0.65 l=0.15
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.1235 ps=1.03 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_1 VPB VNB A1 A2 A3 Y B1 VPWR VGND
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VPB VNB VGND VPWR A1 A2 B1 X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB B1 A1 A2 X B2
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB X A B
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15575 ps=1.355 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_2 VPWR VGND VPB VNB C_N X A B
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_1 VPB VNB VGND VPWR C_N B Y A
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND VPB VNB X A
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_2 VNB VPB VGND VPWR C A Y B
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 X A VPB VNB VGND VPWR
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_4 VNB VPB VGND VPWR A2 A1 B1_N Y
X0 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_33_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.182 ps=1.86 w=0.65 l=0.15
X4 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X11 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B1_N a_33_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X20 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 VPB VNB VGND VPWR B2 A2 A1 B1 X
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 VNB VPB VPWR VGND X A1_N A2_N B2 B1
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.14575 ps=1.335 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20925 pd=1.345 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.20925 ps=1.345 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06615 pd=0.735 as=0.098625 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.098625 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_4 VNB VPB VPWR VGND X S A1 A0
X0 a_204_297# A1 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.16 ps=1.32 w=1 l=0.15
X1 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR S a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_204_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_396_47# A0 a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X6 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.108875 ps=0.985 w=0.65 l=0.15
X7 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_490_47# A1 a_396_47# VNB sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.104 ps=0.97 w=0.65 l=0.15
X11 VGND S a_490_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.274625 ps=1.495 w=0.65 l=0.15
X12 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_396_47# A0 a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.26 ps=1.45 w=0.65 l=0.15
X14 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VPWR S a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X16 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND S a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.108875 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2ai_1 VPB VNB VGND VPWR B1 B2 Y A2_N A1_N
X0 VPWR A2_N a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=1.84 as=0.135 ps=1.27 w=1 l=0.15
X1 Y a_112_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.42 ps=1.84 w=1 l=0.15
X2 VGND B2 a_394_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_112_297# A2_N a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2405 pd=2.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X4 a_112_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17875 ps=1.85 w=0.65 l=0.15
X5 a_112_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X6 VPWR B1 a_478_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X7 a_394_47# a_112_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_394_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_478_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_6 VPB VNB VPWR VGND Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.247 ps=2.06 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.43 ps=2.86 w=1 l=0.15
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VPB VNB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15075 ps=1.345 w=1 l=0.15
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15075 pd=1.345 as=0.074375 ps=0.815 w=0.42 l=0.15
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1304 ps=1.105 w=0.65 l=0.15
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1304 pd=1.105 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 VPB VNB VGND VPWR C B A Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR VPB VNB B C_N A X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_1 VPB VGND VPWR VNB B1 X D1 A1 A2 C1
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.082875 ps=0.905 w=0.65 l=0.15
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.10075 ps=0.96 w=0.65 l=0.15
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.274625 pd=1.495 as=0.2145 ps=1.96 w=0.65 l=0.15
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.082875 pd=0.905 as=0.18525 ps=1.22 w=0.65 l=0.15
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.274625 ps=1.495 w=0.65 l=0.15
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311ai_2 VGND VPWR VPB VNB Y B1 C1 A1 A2 A3
X0 VPWR A1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_55_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y C1 a_729_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.205 ps=1.41 w=1 l=0.15
X4 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_55_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.23075 ps=1.36 w=0.65 l=0.15
X6 VGND A1 a_55_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 a_55_47# B1 a_729_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VGND A2 a_55_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.305 ps=1.61 w=1 l=0.15
X10 VGND A3 a_55_47# VNB sky130_fd_pr__nfet_01v8 ad=0.23075 pd=1.36 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_729_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X12 a_51_297# A2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 a_729_47# B1 a_55_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_301_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_55_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X17 a_51_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y A3 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_301_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_1 VNB VPB VGND VPWR C1 B1 A1 A2 A3 X
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.134875 ps=1.065 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.112125 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125125 ps=1.035 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.134875 pd=1.065 as=0.105625 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.1625 ps=1.325 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1425 ps=1.285 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt clock_divider clk_in clk_out nrst scale[0] scale[1] scale[2] scale[3] scale[4]
+ scale[5] scale[6] scale[7] VPWR VGND
XFILLER_0_7_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0985_ true_scale\[9\] net24 _0004_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_19_Left_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0770_ VGND VPWR _0317_ _0294_ _0292_ _0315_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0968_ VPWR VGND VGND VPWR count\[28\] _0482_ _0481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0899_ VGND VPWR _0436_ count\[5\] count\[4\] _0415_ VPWR VGND sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_4_Left_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0822_ VPWR VGND VGND VPWR true_scale\[23\] _0364_ _0071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0684_ VGND VPWR _0234_ _0236_ _0212_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0753_ VGND VPWR _0299_ _0301_ _0147_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1021_ count\[18\] net27 _0040_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0805_ VPWR VGND VPWR VGND _0348_ _0349_ net21 _0350_ sky130_fd_sc_hd__or3_1
X_0667_ VPWR VGND VGND VPWR _0219_ _0218_ _0220_ sky130_fd_sc_hd__nand2b_1
X_0598_ VGND VPWR _0153_ _0154_ _0129_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0736_ VPWR VGND _0285_ _0284_ _0283_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_38_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0521_ VPWR VGND VPWR VGND net20 net18 net4 _0082_ sky130_fd_sc_hd__or3_4
XFILLER_0_21_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1004_ count\[1\] net23 _0023_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0719_ VPWR VGND VPWR VGND _0241_ _0240_ _0268_ _0269_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_33_Left_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0504_ VPWR VGND VPWR VGND true_scale\[19\] _0068_ true_scale\[18\] _0069_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0984_ true_scale\[8\] net25 _0003_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_20_Left_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0967_ _0481_ net12 _0049_ _0480_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0898_ VGND VPWR _0026_ _0434_ net11 _0435_ VPWR VGND sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_12_Right_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_37_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_30_Right_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0821_ VGND VPWR _0362_ _0363_ count\[23\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0752_ VPWR VGND VGND VPWR _0147_ _0300_ _0299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0683_ VPWR VGND _0235_ _0234_ _0212_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_19_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_129 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1020_ count\[17\] net27 _0039_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0735_ VGND VPWR VPWR VGND _0261_ _0262_ _0284_ _0147_ sky130_fd_sc_hd__a21boi_2
X_0804_ VGND VPWR _0349_ _0340_ _0334_ _0347_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0666_ VPWR VGND VPWR VGND _0196_ _0219_ _0195_ _0197_ sky130_fd_sc_hd__a21boi_1
X_0597_ VGND VPWR VPWR VGND _0150_ _0153_ _0151_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_143 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0520_ VPWR VGND VGND VPWR _0081_ net19 net18 sky130_fd_sc_hd__or2_1
X_1003_ count\[0\] net23 _0022_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_29_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0718_ VPWR VGND VPWR VGND _0249_ _0251_ _0239_ _0268_ sky130_fd_sc_hd__or3_1
X_0649_ VPWR VGND _0203_ _0202_ _0201_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0503_ VPWR VGND VPWR VGND true_scale\[16\] _0066_ true_scale\[17\] true_scale\[15\]
+ _0068_ sky130_fd_sc_hd__or4_2
XFILLER_0_17_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0983_ true_scale\[7\] net23 _0002_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0966_ VGND VPWR _0481_ count\[27\] count\[26\] _0476_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0897_ VPWR VGND VGND VPWR _0435_ count\[4\] _0415_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0820_ VGND VPWR VPWR VGND true_scale\[24\] _0362_ _0072_ sky130_fd_sc_hd__xor2_1
X_0751_ VGND VPWR _0297_ _0299_ _0296_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0682_ VGND VPWR VPWR VGND _0231_ _0234_ _0232_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_34_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0949_ _0468_ _0469_ _0043_ net12 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_33_196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0665_ VPWR VGND _0218_ _0217_ _0214_ VPWR VGND sky130_fd_sc_hd__xor2_2
XFILLER_0_21_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0734_ VGND VPWR _0282_ _0283_ _0147_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0803_ VPWR VGND VPWR VGND _0340_ _0334_ _0347_ _0348_ sky130_fd_sc_hd__a21oi_1
X_0596_ VPWR VGND VGND VPWR _0150_ _0152_ _0151_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_211 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1002_ true_scale\[26\] net29 _0021_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0648_ VGND VPWR _0199_ _0200_ _0202_ _0198_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0717_ VGND VPWR VPWR VGND _0263_ _0267_ _0264_ sky130_fd_sc_hd__xor2_1
X_0579_ VGND VPWR _0135_ _0136_ _0129_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_203 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0502_ VPWR VGND VGND VPWR true_scale\[15\] _0066_ _0067_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_84 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0982_ true_scale\[6\] net25 _0001_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0965_ VPWR VGND VGND VPWR _0480_ count\[27\] _0478_ sky130_fd_sc_hd__or2_1
X_0896_ VPWR VGND VGND VPWR count\[4\] _0434_ _0415_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0681_ VPWR VGND _0233_ _0232_ _0231_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0750_ VPWR VGND VGND VPWR _0297_ _0296_ _0298_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_19_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0948_ VPWR VGND VGND VPWR _0469_ count\[21\] _0466_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0879_ VPWR VGND VPWR VGND _0402_ _0420_ _0404_ _0401_ _0421_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0802_ _0347_ _0345_ _0346_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_0664_ VGND VPWR _0217_ _0094_ _0215_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_76 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0733_ VGND VPWR VPWR VGND _0279_ _0282_ _0280_ sky130_fd_sc_hd__xor2_1
X_0595_ VGND VPWR VPWR VGND _0151_ net18 net20 _0057_ _0095_ _0130_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1001_ true_scale\[25\] net28 _0020_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0647_ VPWR VGND VPWR VGND _0199_ _0200_ _0198_ _0201_ sky130_fd_sc_hd__or3_1
X_0578_ VGND VPWR _0133_ _0135_ _0131_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0716_ VPWR VGND VPWR VGND _0266_ _0265_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0501_ VPWR VGND VPWR VGND true_scale\[13\] _0064_ true_scale\[14\] true_scale\[12\]
+ _0066_ sky130_fd_sc_hd__or4_2
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0981_ true_scale\[5\] net25 _0000_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0964_ _0478_ _0479_ _0048_ net12 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0895_ _0415_ net11 _0025_ _0433_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0680_ VPWR VGND VPWR VGND _0217_ _0214_ _0216_ _0232_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_24_Left_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0947_ VPWR VGND _0468_ _0466_ count\[21\] VPWR VGND sky130_fd_sc_hd__and2_1
X_0878_ VPWR VGND VPWR VGND _0407_ _0419_ _0406_ _0420_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0801_ VPWR VGND VGND VPWR _0328_ _0346_ _0344_ _0343_ _0330_ sky130_fd_sc_hd__o211ai_1
X_0663_ _0216_ _0215_ _0094_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_0594_ VGND VPWR VPWR VGND _0080_ _0150_ _0148_ sky130_fd_sc_hd__xor2_1
X_0732_ VPWR VGND _0281_ _0280_ _0279_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_15_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1000_ true_scale\[24\] net28 _0019_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_54 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0715_ VPWR VGND VGND VPWR _0265_ _0263_ _0264_ sky130_fd_sc_hd__or2_1
X_0646_ VPWR VGND VPWR VGND _0178_ _0172_ _0177_ _0200_ sky130_fd_sc_hd__a21oi_1
X_0577_ _0134_ _0133_ _0131_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_11_Left_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0500_ VPWR VGND VGND VPWR true_scale\[12\] _0064_ _0065_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_28_Right_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0629_ VGND VPWR _0183_ _0184_ _0147_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0980_ VPWR VGND VPWR VGND _0429_ _0055_ _0489_ _0054_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0894_ VPWR VGND _0433_ count\[2\] count\[1\] count\[0\] count\[3\] VGND VPWR sky130_fd_sc_hd__a31o_1
X_0963_ VPWR VGND VGND VPWR _0479_ count\[26\] _0476_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0877_ VPWR VGND VPWR VGND _0410_ _0412_ _0409_ _0419_ _0418_ sky130_fd_sc_hd__or4b_1
X_0946_ _0466_ _0467_ _0042_ net12 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_41_Left_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_18_163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0800_ VPWR VGND VPWR VGND _0345_ _0330_ _0328_ _0343_ _0344_ sky130_fd_sc_hd__a211oi_1
X_0731_ VPWR VGND VPWR VGND _0258_ _0128_ _0257_ _0280_ sky130_fd_sc_hd__a21o_1
X_0662_ VGND VPWR _0215_ _0090_ _0096_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_0593_ _0149_ _0077_ _0078_ _0079_ _0148_ VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_0929_ _0456_ count\[15\] count\[13\] count\[14\] _0450_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
XFILLER_0_15_188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_32_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0645_ VPWR VGND VPWR VGND _0197_ _0196_ _0195_ _0199_ sky130_fd_sc_hd__a21oi_1
X_0714_ VGND VPWR VPWR VGND _0246_ _0264_ net9 _0111_ _0247_ sky130_fd_sc_hd__a31oi_2
X_0576_ VGND VPWR VGND VPWR _0115_ _0095_ _0133_ _0132_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0628_ VGND VPWR VPWR VGND _0180_ _0183_ _0181_ sky130_fd_sc_hd__xor2_1
X_0559_ VGND VPWR _0081_ _0095_ _0117_ _0097_ VPWR VGND sky130_fd_sc_hd__o21ai_2
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0962_ VPWR VGND _0478_ _0476_ count\[26\] VPWR VGND sky130_fd_sc_hd__and2_1
X_0893_ VGND VPWR _0024_ net11 _0414_ _0432_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_36_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_19_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0876_ VGND VPWR _0418_ _0416_ _0415_ _0417_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0945_ VPWR VGND VPWR VGND _0462_ count\[19\] count\[20\] _0467_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_175 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_33_178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_112 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0730_ VGND VPWR _0278_ _0279_ _0128_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0661_ VPWR VGND VGND VPWR _0212_ _0213_ _0214_ sky130_fd_sc_hd__nor2_1
X_0592_ VPWR VGND _0148_ net17 net7 VPWR VGND sky130_fd_sc_hd__xor2_2
X_0928_ _0454_ _0455_ _0036_ net13 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0859_ VGND VPWR _0401_ _0063_ count\[9\] _0400_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_30_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0644_ VGND VPWR _0198_ _0196_ _0195_ _0197_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_12_115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0713_ VGND VPWR _0262_ _0263_ _0147_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0575_ VGND VPWR _0132_ _0058_ net19 net18 VPWR VGND sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_1_Right_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_210 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_7_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0627_ VPWR VGND _0182_ _0181_ _0180_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0558_ VGND VPWR _0116_ _0095_ _0115_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0961_ _0476_ _0477_ _0047_ net12 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0892_ VPWR VGND VPWR VGND count\[1\] count\[0\] count\[2\] _0432_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0944_ VGND VPWR _0466_ count\[20\] count\[19\] _0462_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ VPWR VGND VGND VPWR count\[4\] _0417_ true_scale\[5\] sky130_fd_sc_hd__nand2_1
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0591_ VGND VPWR VPWR VGND _0112_ _0147_ _0060_ _0114_ sky130_fd_sc_hd__o21ai_4
X_0660_ VPWR VGND VGND VPWR net10 _0084_ _0213_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ VPWR VGND VPWR VGND _0450_ count\[13\] count\[14\] _0455_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0789_ VPWR VGND VGND VPWR _0332_ _0333_ _0335_ sky130_fd_sc_hd__nand2b_1
X_0858_ VGND VPWR _0062_ true_scale\[10\] _0400_ true_scale\[9\] VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0643_ VGND VPWR VGND VPWR _0197_ _0175_ _0093_ _0091_ _0089_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_12_127 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0574_ VGND VPWR _0130_ _0131_ _0096_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0712_ VGND VPWR VPWR VGND _0259_ _0262_ _0260_ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_230 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0626_ VGND VPWR VGND VPWR _0181_ _0153_ _0128_ _0152_ sky130_fd_sc_hd__a21bo_1
X_0557_ VGND VPWR VPWR VGND _0079_ _0088_ _0078_ _0115_ sky130_fd_sc_hd__or3_2
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0609_ VGND VPWR _0165_ _0163_ _0142_ _0164_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0960_ VPWR VGND VGND VPWR _0477_ count\[25\] _0474_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0891_ VGND VPWR _0023_ net11 _0413_ _0431_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_14_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_36_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_36_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0874_ VPWR VGND VGND VPWR _0416_ count\[4\] true_scale\[5\] sky130_fd_sc_hd__or2_1
X_0943_ VGND VPWR _0041_ _0464_ net13 _0465_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_27_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Left_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0590_ VGND VPWR VPWR VGND _0007_ _0146_ net16 true_scale\[12\] sky130_fd_sc_hd__mux2_1
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0926_ VGND VPWR _0454_ count\[14\] count\[13\] _0450_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0857_ VGND VPWR VPWR VGND count\[10\] _0399_ _0398_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0788_ VPWR VGND VGND VPWR _0333_ _0332_ _0334_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0711_ VPWR VGND VGND VPWR _0259_ _0261_ _0260_ sky130_fd_sc_hd__nand2_1
X_0642_ VGND VPWR VGND VPWR _0196_ _0175_ _0093_ _0089_ _0091_ sky130_fd_sc_hd__a211o_1
X_0573_ VPWR VGND VPWR VGND _0075_ _0130_ _0081_ _0097_ sky130_fd_sc_hd__a21boi_1
X_0909_ VPWR VGND VPWR VGND _0438_ count\[7\] count\[8\] _0443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0625_ VGND VPWR _0179_ _0180_ _0172_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0556_ VPWR VGND VPWR VGND _0114_ _0113_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0608_ VPWR VGND VGND VPWR _0108_ _0164_ _0128_ sky130_fd_sc_hd__nand2_1
X_0539_ VGND VPWR VGND VPWR _0097_ net19 net18 _0098_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_24_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ VPWR VGND VGND VPWR _0431_ count\[0\] count\[1\] sky130_fd_sc_hd__or2_1
XFILLER_0_36_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0873_ _0415_ count\[3\] count\[0\] count\[1\] count\[2\] VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_0942_ VPWR VGND VGND VPWR _0465_ count\[19\] _0462_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_33_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_24_104 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_24_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0787_ VPWR VGND VPWR VGND _0319_ _0191_ _0316_ _0333_ sky130_fd_sc_hd__a21oi_1
X_0925_ VGND VPWR _0035_ _0452_ net13 _0453_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0856_ VGND VPWR _0063_ _0398_ true_scale\[11\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0641_ VGND VPWR _0195_ _0060_ _0194_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_0710_ VPWR VGND VPWR VGND _0119_ _0118_ _0260_ _0129_ sky130_fd_sc_hd__o21bai_1
X_0572_ VGND VPWR VGND VPWR _0129_ _0113_ net10 sky130_fd_sc_hd__xnor2_4
XFILLER_0_7_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0908_ VGND VPWR _0442_ count\[8\] count\[7\] _0438_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0839_ VGND VPWR _0380_ _0381_ count\[17\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_210 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0624_ VPWR VGND VGND VPWR _0177_ _0178_ _0179_ sky130_fd_sc_hd__nand2b_1
X_0555_ VGND VPWR VGND VPWR _0111_ _0113_ net9 sky130_fd_sc_hd__xor2_4
XPHY_EDGE_ROW_5_Right_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0607_ VPWR VGND VPWR VGND _0121_ _0122_ _0105_ _0163_ _0141_ sky130_fd_sc_hd__or4b_1
X_0538_ VGND VPWR VPWR VGND net20 net18 _0097_ net19 sky130_fd_sc_hd__a21boi_2
XFILLER_0_39_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout20 VPWR VGND net20 net3 VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0941_ VPWR VGND VGND VPWR count\[19\] _0464_ _0462_ sky130_fd_sc_hd__nand2_1
X_0872_ VPWR VGND VGND VPWR count\[0\] count\[1\] _0414_ count\[2\] sky130_fd_sc_hd__nand3_1
XFILLER_0_41_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_24_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0924_ VPWR VGND VGND VPWR _0453_ count\[13\] _0450_ sky130_fd_sc_hd__or2_1
X_0786_ VPWR VGND VGND VPWR _0330_ _0331_ _0332_ sky130_fd_sc_hd__nor2_1
X_0855_ VGND VPWR _0396_ _0397_ count\[11\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0640_ VPWR VGND VGND VPWR _0192_ _0193_ _0194_ sky130_fd_sc_hd__nor2_1
X_0571_ VGND VPWR VGND VPWR _0128_ _0113_ _0060_ sky130_fd_sc_hd__xnor2_4
X_0907_ VGND VPWR _0029_ _0440_ net11 _0441_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0769_ VPWR VGND VPWR VGND _0294_ _0292_ _0315_ _0316_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0838_ VGND VPWR VPWR VGND true_scale\[18\] _0380_ _0068_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0554_ VPWR VGND VGND VPWR _0112_ net9 _0111_ sky130_fd_sc_hd__nand2_2
X_0623_ VGND VPWR VGND VPWR _0178_ _0176_ _0088_ _0175_ _0149_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0537_ VGND VPWR VGND VPWR _0096_ _0086_ net17 sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0606_ VPWR VGND VPWR VGND _0140_ _0138_ _0159_ _0162_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_49 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout21 VPWR VGND net21 net22 VPWR VGND sky130_fd_sc_hd__buf_2
X_0940_ _0462_ _0463_ _0040_ net13 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0871_ VPWR VGND VGND VPWR count\[0\] _0413_ count\[1\] sky130_fd_sc_hd__nand2_1
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0923_ VPWR VGND VGND VPWR count\[13\] _0452_ _0450_ sky130_fd_sc_hd__nand2_1
X_0854_ VPWR VGND VGND VPWR _0065_ _0395_ _0396_ sky130_fd_sc_hd__nor2_1
X_0785_ _0331_ _0211_ _0329_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_0_36_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_21_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0570_ VGND VPWR VPWR VGND _0006_ _0127_ net16 true_scale\[11\] sky130_fd_sc_hd__mux2_1
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_28_220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0906_ VPWR VGND VGND VPWR _0441_ count\[7\] _0438_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0837_ VPWR VGND VGND VPWR _0379_ _0377_ _0378_ sky130_fd_sc_hd__or2_1
X_0768_ VGND VPWR _0195_ _0315_ net7 VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0699_ VGND VPWR _0235_ _0248_ _0250_ _0233_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_0622_ VGND VPWR VGND VPWR _0177_ _0088_ _0149_ _0175_ _0176_ sky130_fd_sc_hd__o211a_1
X_0553_ VGND VPWR VGND VPWR _0086_ net17 _0084_ _0111_ sky130_fd_sc_hd__a21o_2
XFILLER_0_17_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0605_ VPWR VGND VPWR VGND _0140_ _0138_ _0159_ _0161_ sky130_fd_sc_hd__a21oi_1
X_0536_ VGND VPWR VGND VPWR _0086_ _0095_ net17 sky130_fd_sc_hd__xor2_4
X_1019_ count\[16\] net27 _0038_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_30_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0519_ VGND VPWR VPWR VGND _0002_ _0080_ net16 true_scale\[7\] sky130_fd_sc_hd__mux2_1
Xfanout11 VGND VPWR net14 net11 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout22 VGND VPWR net2 net22 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ VGND VPWR _0411_ _0412_ count\[5\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0999_ true_scale\[23\] net28 _0018_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Left_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0922_ _0450_ _0451_ _0034_ net14 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0853_ VPWR VGND _0395_ _0064_ true_scale\[12\] VPWR VGND sky130_fd_sc_hd__and2_1
X_0784_ _0330_ _0329_ _0211_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
Xinput1 VGND VPWR net1 clk_in VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_37_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0905_ VPWR VGND VGND VPWR count\[7\] _0440_ _0438_ sky130_fd_sc_hd__nand2_1
X_0836_ VPWR VGND VPWR VGND _0376_ _0069_ count\[18\] _0378_ sky130_fd_sc_hd__a21oi_1
X_0767_ VPWR VGND net21 _0312_ _0313_ _0016_ _0314_ VPWR VGND sky130_fd_sc_hd__o31ai_1
X_0698_ VPWR VGND VGND VPWR _0233_ _0235_ _0248_ _0249_ sky130_fd_sc_hd__o21a_1
X_0621_ VGND VPWR VGND VPWR _0176_ _0089_ _0082_ _0174_ sky130_fd_sc_hd__a21bo_1
X_0552_ VPWR VGND VPWR VGND _0109_ true_scale\[10\] net22 _0005_ _0110_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1035_ signal_clk_out net29 _0054_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_10_Left_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0819_ VGND VPWR VPWR VGND true_scale\[26\] _0361_ _0073_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_9_Right_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0604_ VGND VPWR _0160_ _0140_ _0138_ _0159_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0535_ VPWR VGND VPWR VGND _0094_ _0088_ _0093_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1018_ count\[15\] net27 _0037_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_30_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0518_ VPWR VGND VPWR VGND _0078_ _0079_ _0077_ _0080_ sky130_fd_sc_hd__or3_1
Xfanout23 VGND VPWR net24 net23 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout12 VGND VPWR net13 net12 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0998_ true_scale\[22\] net28 _0017_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_174 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0921_ VPWR VGND VGND VPWR _0451_ count\[12\] _0448_ sky130_fd_sc_hd__or2_1
X_0783_ VPWR VGND VGND VPWR _0329_ _0327_ _0328_ sky130_fd_sc_hd__or2_1
X_0852_ VGND VPWR _0393_ _0394_ count\[12\] VPWR VGND sky130_fd_sc_hd__xnor2_1
Xinput2 VGND VPWR net2 nrst VPWR VGND sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_40_Left_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_200 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_20_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0904_ _0438_ _0439_ _0028_ net11 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_52 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0835_ VGND VPWR _0377_ _0069_ count\[18\] _0376_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0766_ VPWR VGND VGND VPWR true_scale\[21\] _0314_ net21 sky130_fd_sc_hd__nand2_1
X_0697_ VGND VPWR _0247_ _0248_ _0112_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0620_ VPWR VGND VPWR VGND _0082_ _0175_ _0174_ _0088_ sky130_fd_sc_hd__or3b_2
X_0551_ VPWR VGND VPWR VGND _0107_ _0106_ net22 _0110_ sky130_fd_sc_hd__a21oi_1
X_1034_ count\[31\] net26 _0053_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0818_ VPWR VGND VPWR VGND _0356_ _0073_ count\[24\] _0360_ sky130_fd_sc_hd__a21oi_1
X_0749_ VPWR VGND VGND VPWR _0129_ _0278_ _0277_ _0297_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0534_ VGND VPWR _0093_ _0086_ _0082_ _0089_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0603_ VGND VPWR _0157_ _0159_ _0147_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_222 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_1017_ count\[14\] net27 _0036_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0517_ _0079_ net18 net20 VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
Xfanout24 VGND VPWR net25 net24 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout13 VGND VPWR net14 net13 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0997_ true_scale\[21\] net28 _0016_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0920_ _0450_ count\[12\] count\[10\] count\[11\] _0444_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_0782_ VGND VPWR _0328_ _0195_ net7 _0326_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0851_ VGND VPWR _0065_ _0393_ true_scale\[13\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Right_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xinput3 VGND VPWR net3 scale[0] VPWR VGND sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_27_Right_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_14_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_14_153 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0903_ VPWR VGND VGND VPWR _0439_ count\[6\] _0436_ sky130_fd_sc_hd__or2_1
X_0834_ VGND VPWR _0068_ true_scale\[19\] _0376_ true_scale\[18\] VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0765_ VPWR VGND VGND VPWR _0305_ _0311_ _0313_ sky130_fd_sc_hd__nor2_1
X_0696_ VGND VPWR VPWR VGND _0244_ _0247_ _0245_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0550_ VPWR VGND VPWR VGND _0109_ _0108_ sky130_fd_sc_hd__inv_2
X_1033_ count\[30\] net26 _0052_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0817_ VPWR VGND _0359_ _0358_ count\[31\] count\[26\] _0074_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0748_ VPWR VGND _0296_ _0295_ _0294_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0679_ VGND VPWR _0230_ _0231_ _0113_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_0_Right_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0533_ VPWR VGND VPWR VGND _0089_ _0085_ _0091_ _0092_ sky130_fd_sc_hd__a21o_1
X_0602_ VPWR VGND VGND VPWR _0147_ _0158_ _0157_ sky130_fd_sc_hd__nand2_1
X_1016_ count\[13\] net27 _0035_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_148 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0516_ VPWR VGND VGND VPWR net18 net20 _0078_ net19 sky130_fd_sc_hd__nor3b_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xfanout25 VPWR VGND VPWR VGND net25 net1 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout14 VGND VPWR _0430_ net14 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0996_ true_scale\[20\] net28 _0015_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ VGND VPWR VPWR VGND count\[13\] _0392_ _0391_ sky130_fd_sc_hd__xor2_1
X_0781_ VPWR VGND VPWR VGND _0195_ net7 _0326_ _0327_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_23_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 VGND VPWR net4 scale[1] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0979_ VGND VPWR _0429_ net22 _0489_ _0055_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_27_Left_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0902_ _0438_ count\[6\] count\[4\] count\[5\] _0415_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_0833_ VPWR VGND VGND VPWR _0375_ _0373_ _0374_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0764_ VPWR VGND _0312_ _0311_ _0305_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0695_ VPWR VGND _0246_ _0245_ _0244_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1032_ count\[29\] net26 _0051_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0816_ _0358_ count\[29\] count\[27\] count\[28\] count\[30\] VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_1
X_0747_ VPWR VGND VGND VPWR _0173_ _0295_ _0293_ sky130_fd_sc_hd__nand2_1
X_0678_ VGND VPWR VGND VPWR _0230_ _0229_ _0100_ _0099_ sky130_fd_sc_hd__a21bo_1
X_0601_ VGND VPWR _0155_ _0157_ _0154_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0532_ VPWR VGND VPWR VGND _0089_ _0082_ _0086_ _0091_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ count\[12\] net25 _0034_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_14_Left_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0515_ _0077_ net18 net19 VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
Xfanout26 VGND VPWR net27 net26 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout15 VPWR VGND net15 net16 VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_0_25_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0995_ true_scale\[19\] net28 _0014_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_188 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_17_196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0780_ VGND VPWR VPWR VGND net17 _0326_ net10 sky130_fd_sc_hd__xor2_1
XFILLER_0_11_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_23_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 VGND VPWR net5 scale[2] VPWR VGND sky130_fd_sc_hd__buf_1
XFILLER_0_36_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0978_ VGND VPWR _0053_ _0487_ net12 _0488_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0901_ _0436_ _0437_ _0027_ net11 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_11_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0832_ VPWR VGND VPWR VGND _0372_ _0070_ count\[19\] _0374_ sky130_fd_sc_hd__a21oi_1
X_0763_ VPWR VGND VPWR VGND _0309_ _0310_ _0308_ _0311_ sky130_fd_sc_hd__or3_1
X_0694_ VPWR VGND VPWR VGND _0229_ _0099_ _0113_ _0245_ _0100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_19_236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_1031_ count\[28\] net26 _0050_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0746_ VPWR VGND VGND VPWR _0294_ _0173_ _0293_ sky130_fd_sc_hd__or2_1
X_0815_ VGND VPWR VPWR VGND _0357_ _0356_ _0073_ count\[24\] _0355_ _0074_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0677_ VPWR VGND VPWR VGND _0095_ _0082_ _0088_ _0229_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0531_ VPWR VGND VGND VPWR _0082_ _0090_ _0089_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0600_ VPWR VGND VGND VPWR _0155_ _0154_ _0156_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1014_ count\[11\] net24 _0033_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0729_ VGND VPWR _0276_ _0278_ _0275_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_31_Left_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0514_ VPWR VGND VPWR VGND _0075_ true_scale\[6\] net22 _0001_ _0076_ sky130_fd_sc_hd__a22o_1
Xfanout27 VPWR VGND net27 net29 VPWR VGND sky130_fd_sc_hd__buf_2
Xfanout16 VGND VPWR _0056_ net16 VPWR VGND sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_44 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0994_ true_scale\[18\] net28 _0013_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 VGND VPWR scale[3] net6 VPWR VGND sky130_fd_sc_hd__clkbuf_4
X_0977_ VPWR VGND VGND VPWR count\[31\] _0488_ _0486_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_14_Right_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_20_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0900_ VPWR VGND VPWR VGND _0415_ count\[4\] count\[5\] _0437_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_32_Right_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_11_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0831_ VGND VPWR _0373_ _0070_ count\[19\] _0372_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0762_ VGND VPWR VGND VPWR _0285_ _0266_ _0286_ _0310_ sky130_fd_sc_hd__o21ba_1
X_0693_ VGND VPWR _0128_ _0244_ _0119_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_41_Right_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1030_ count\[27\] net26 _0049_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0814_ VGND VPWR _0072_ true_scale\[25\] _0356_ true_scale\[24\] VPWR VGND sky130_fd_sc_hd__o21ai_1
X_0676_ VPWR VGND VGND VPWR true_scale\[16\] net15 _0228_ _0011_ sky130_fd_sc_hd__o21a_1
X_0745_ VPWR VGND VGND VPWR _0291_ _0293_ _0292_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_232 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0530_ VGND VPWR VGND VPWR net5 net4 _0089_ net3 sky130_fd_sc_hd__nand3_2
XFILLER_0_0_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1013_ count\[10\] net24 _0032_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_4_Right_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0728_ VPWR VGND VGND VPWR _0277_ _0275_ _0276_ sky130_fd_sc_hd__or2_1
X_0659_ VPWR VGND VGND VPWR _0060_ _0085_ _0212_ sky130_fd_sc_hd__nor2_1
X_0513_ VPWR VGND VPWR VGND net20 net19 net22 _0076_ sky130_fd_sc_hd__a21oi_1
Xfanout17 net17 net8 VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout28 VGND VPWR net29 net28 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0993_ true_scale\[17\] net27 _0012_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 VPWR VGND net7 scale[4] VPWR VGND sky130_fd_sc_hd__buf_4
X_0976_ VPWR VGND VGND VPWR _0487_ count\[31\] _0486_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_238 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_9_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0830_ VPWR VGND VGND VPWR true_scale\[20\] _0372_ _0069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0692_ VGND VPWR VPWR VGND _0012_ _0243_ net15 true_scale\[17\] sky130_fd_sc_hd__mux2_1
X_0761_ VGND VPWR _0309_ _0270_ _0267_ _0288_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_12_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0959_ VGND VPWR _0476_ count\[25\] count\[24\] _0472_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_10_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xinput10 VPWR VGND net10 scale[7] VPWR VGND sky130_fd_sc_hd__buf_4
X_0813_ VPWR VGND VPWR VGND count\[27\] _0354_ count\[26\] _0355_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0744_ VPWR VGND VGND VPWR _0292_ _0174_ _0273_ sky130_fd_sc_hd__or2_1
X_0675_ VGND VPWR _0227_ net15 _0228_ _0226_ VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_241 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_1012_ count\[9\] net24 _0031_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0727_ VPWR VGND VPWR VGND _0255_ _0095_ _0088_ _0276_ sky130_fd_sc_hd__a21oi_1
X_0658_ VGND VPWR VGND VPWR _0192_ _0060_ _0193_ _0211_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_40_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0589_ VGND VPWR _0145_ _0146_ _0144_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0512_ VPWR VGND VGND VPWR _0075_ net19 net20 sky130_fd_sc_hd__or2_1
Xfanout18 VGND VPWR net5 net18 VPWR VGND sky130_fd_sc_hd__clkbuf_2
Xfanout29 VPWR VGND VPWR VGND net29 net1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_20_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0992_ true_scale\[16\] net27 _0011_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 VGND VPWR net8 scale[5] VPWR VGND sky130_fd_sc_hd__buf_1
X_0975_ _0486_ net12 _0052_ _0485_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_14_103 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0760_ VPWR VGND VPWR VGND _0308_ _0268_ _0307_ _0241_ _0306_ sky130_fd_sc_hd__a211oi_1
X_0691_ VGND VPWR VPWR VGND _0239_ _0243_ _0242_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0889_ _0022_ count\[0\] net11 VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
X_0958_ _0474_ _0475_ _0046_ net13 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_6_Left_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0812_ VPWR VGND VPWR VGND count\[29\] count\[31\] count\[30\] count\[28\] _0354_
+ sky130_fd_sc_hd__or4_1
X_0743_ VPWR VGND VGND VPWR _0174_ _0291_ _0273_ sky130_fd_sc_hd__nand2_1
X_0674_ VPWR VGND VPWR VGND _0208_ _0206_ _0225_ _0227_ sky130_fd_sc_hd__a21oi_1
X_1011_ count\[8\] net23 _0030_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0726_ VPWR VGND VGND VPWR _0273_ _0275_ _0274_ sky130_fd_sc_hd__nand2_1
X_0588_ VPWR VGND VGND VPWR _0109_ _0126_ _0124_ _0145_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0657_ VGND VPWR VGND VPWR _0210_ _0202_ _0191_ _0201_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_9_Left_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0511_ VGND VPWR VPWR VGND _0000_ true_scale\[5\] net22 net20 sky130_fd_sc_hd__mux2_1
Xfanout19 VPWR VGND net19 net4 VPWR VGND sky130_fd_sc_hd__buf_2
X_0709_ VGND VPWR _0258_ _0259_ _0129_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_35_Left_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ true_scale\[15\] net28 _0010_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_181 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xinput9 VPWR VGND net9 scale[6] VPWR VGND sky130_fd_sc_hd__buf_4
XFILLER_0_36_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0974_ VPWR VGND _0486_ _0484_ count\[30\] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_13_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0690_ VPWR VGND _0242_ _0241_ _0240_ VPWR VGND sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_22_Left_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Right_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_6_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0957_ VPWR VGND VGND VPWR _0475_ count\[24\] _0472_ sky130_fd_sc_hd__or2_1
X_0888_ VPWR VGND _0430_ _0429_ net2 VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_10_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0673_ VGND VPWR _0226_ _0208_ _0206_ _0225_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0742_ VPWR VGND VGND VPWR _0290_ net16 true_scale\[20\] _0289_ _0015_ sky130_fd_sc_hd__o22a_1
X_0811_ VGND VPWR VPWR VGND _0021_ _0353_ _0343_ true_scale\[26\] net15 sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1010_ count\[7\] net23 _0029_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_213 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0656_ VPWR VGND _0010_ _0209_ _0208_ net15 _0190_ VGND VPWR sky130_fd_sc_hd__a31o_1
X_0725_ VPWR VGND VGND VPWR _0274_ net5 _0148_ sky130_fd_sc_hd__or2_1
X_0587_ VPWR VGND _0144_ _0143_ _0142_ VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0510_ VGND VPWR VPWR VGND clk_out _0074_ signal_clk_out net28 sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_8_Right_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0639_ VGND VPWR _0193_ net17 net6 net9 VPWR VGND sky130_fd_sc_hd__and3_1
X_0708_ VGND VPWR VPWR VGND _0133_ _0258_ _0256_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0990_ true_scale\[14\] net24 _0009_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0973_ VPWR VGND VGND VPWR _0485_ count\[30\] _0484_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0956_ VPWR VGND _0474_ _0472_ count\[24\] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_27_241 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0887_ VPWR VGND VPWR VGND _0428_ _0360_ _0357_ _0429_ _0359_ sky130_fd_sc_hd__or4b_1
XFILLER_0_10_185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0810_ VPWR VGND VPWR VGND _0352_ true_scale\[25\] net21 _0020_ _0353_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0672_ VGND VPWR _0222_ _0225_ _0210_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0741_ VPWR VGND _0290_ _0288_ _0271_ _0265_ net21 VGND VPWR sky130_fd_sc_hd__a31o_1
X_0939_ VPWR VGND VGND VPWR _0463_ count\[18\] _0460_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_225 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_8_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0586_ VPWR VGND VGND VPWR _0143_ _0121_ _0141_ sky130_fd_sc_hd__or2_1
X_0655_ VPWR VGND VGND VPWR _0188_ _0207_ _0209_ sky130_fd_sc_hd__nand2b_1
X_0724_ VPWR VGND VGND VPWR net5 _0273_ _0148_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_100 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0707_ VPWR VGND VGND VPWR _0133_ _0256_ _0257_ sky130_fd_sc_hd__nor2_1
X_0638_ VGND VPWR VGND VPWR net17 net6 _0192_ net9 sky130_fd_sc_hd__a21oi_2
X_0569_ VGND VPWR _0126_ _0127_ _0108_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_40_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0972_ _0484_ net12 _0051_ _0483_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_37_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0955_ _0472_ _0473_ _0045_ net13 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0886_ VGND VPWR _0361_ _0427_ _0428_ count\[25\] VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0740_ VPWR VGND VPWR VGND _0271_ _0265_ _0288_ _0289_ sky130_fd_sc_hd__a21oi_1
X_0671_ VPWR VGND VGND VPWR _0210_ _0222_ _0224_ sky130_fd_sc_hd__nor2_1
X_0938_ _0462_ count\[18\] count\[16\] count\[17\] _0456_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_0869_ VGND VPWR VPWR VGND true_scale\[5\] _0411_ true_scale\[6\] sky130_fd_sc_hd__xor2_1
XFILLER_0_30_204 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_28_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0723_ VPWR VGND VPWR VGND _0271_ true_scale\[19\] net21 _0014_ _0272_ sky130_fd_sc_hd__a22o_1
X_0585_ VPWR VGND VGND VPWR _0121_ _0142_ _0141_ sky130_fd_sc_hd__nand2_1
X_0654_ VPWR VGND VPWR VGND _0187_ _0185_ _0207_ _0208_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0706_ VGND VPWR _0255_ _0256_ _0095_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0637_ VGND VPWR VGND VPWR _0169_ _0060_ _0170_ _0191_ sky130_fd_sc_hd__o21bai_4
X_0499_ VPWR VGND VPWR VGND true_scale\[10\] _0062_ true_scale\[11\] true_scale\[9\]
+ _0064_ sky130_fd_sc_hd__or4_1
X_0568_ VPWR VGND VGND VPWR _0124_ _0126_ _0125_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_28 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0971_ VGND VPWR _0484_ count\[29\] count\[28\] _0481_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_26_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0954_ VPWR VGND _0473_ _0466_ count\[22\] count\[21\] count\[23\] VGND VPWR sky130_fd_sc_hd__a31o_1
X_0885_ VPWR VGND VPWR VGND _0427_ _0426_ _0363_ count\[25\] _0361_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0670_ VPWR VGND VGND VPWR _0210_ _0223_ _0222_ sky130_fd_sc_hd__nand2_1
X_0799_ VPWR VGND VPWR VGND net10 net8 net9 _0344_ sky130_fd_sc_hd__a21o_1
X_0937_ _0460_ _0461_ _0039_ net13 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0868_ VPWR VGND VPWR VGND _0408_ _0061_ count\[6\] _0410_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_238 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0653_ VGND VPWR _0207_ _0204_ _0205_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_0722_ _0272_ _0267_ _0269_ _0270_ net16 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
X_0584_ VGND VPWR _0139_ _0141_ _0112_ VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0636_ VPWR VGND _0190_ net21 true_scale\[15\] VPWR VGND sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_29_Left_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0705_ VPWR VGND VPWR VGND _0081_ net19 _0058_ _0255_ _0097_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_13_Left_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0498_ VPWR VGND VPWR VGND true_scale\[10\] _0062_ true_scale\[9\] _0063_ sky130_fd_sc_hd__or3_1
X_0567_ VPWR VGND VGND VPWR _0105_ _0125_ _0123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_41_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0619_ VGND VPWR net17 _0174_ net6 VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0970_ VPWR VGND VPWR VGND _0481_ count\[28\] count\[29\] _0483_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0953_ VGND VPWR _0472_ count\[23\] count\[22\] _0468_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0884_ VPWR VGND VPWR VGND _0366_ _0425_ _0369_ _0365_ _0426_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0936_ VPWR VGND VPWR VGND _0456_ count\[16\] count\[17\] _0461_ sky130_fd_sc_hd__a21o_1
X_0798_ VPWR VGND VGND VPWR net8 net9 _0343_ net10 sky130_fd_sc_hd__nand3_1
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0867_ VGND VPWR _0409_ _0061_ count\[6\] _0408_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_12_239 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0583_ VPWR VGND VGND VPWR _0112_ _0139_ _0140_ sky130_fd_sc_hd__nand2b_1
X_0652_ VPWR VGND VGND VPWR _0206_ _0204_ _0205_ sky130_fd_sc_hd__or2_1
X_0721_ VGND VPWR _0270_ _0267_ _0271_ _0269_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_0919_ _0448_ _0449_ _0033_ net14 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_0_29_147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_20_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0566_ VPWR VGND VGND VPWR _0124_ _0105_ _0123_ sky130_fd_sc_hd__or2_1
X_0635_ VPWR VGND VGND VPWR _0188_ _0189_ _0009_ net22 true_scale\[14\] sky130_fd_sc_hd__o2bb2ai_1
X_0704_ VGND VPWR VPWR VGND _0013_ _0254_ net15 true_scale\[18\] sky130_fd_sc_hd__mux2_1
X_0497_ VPWR VGND VPWR VGND true_scale\[6\] true_scale\[8\] true_scale\[7\] true_scale\[5\]
+ _0062_ sky130_fd_sc_hd__or4_2
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0618_ VGND VPWR _0171_ _0173_ _0060_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0549_ VPWR VGND VGND VPWR _0106_ _0107_ _0108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_39_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0952_ VGND VPWR _0044_ _0470_ net12 _0471_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0883_ VPWR VGND VPWR VGND _0375_ _0424_ _0379_ _0371_ _0425_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_33_215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0935_ VGND VPWR _0460_ count\[17\] count\[16\] _0456_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0866_ VGND VPWR true_scale\[6\] true_scale\[7\] _0408_ true_scale\[5\] VPWR VGND
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0797_ VPWR VGND _0018_ _0341_ _0340_ net15 _0342_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_3_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0720_ VPWR VGND VPWR VGND _0250_ _0238_ _0251_ _0270_ sky130_fd_sc_hd__a21oi_1
X_0582_ VGND VPWR _0137_ _0139_ _0136_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0651_ VPWR VGND VPWR VGND _0183_ _0147_ _0182_ _0205_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0918_ VPWR VGND VPWR VGND _0444_ count\[10\] count\[11\] _0449_ sky130_fd_sc_hd__a21o_1
X_0849_ VPWR VGND VGND VPWR _0066_ _0391_ _0390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0703_ VGND VPWR _0253_ _0254_ _0252_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0496_ VPWR VGND VPWR VGND true_scale\[6\] true_scale\[7\] true_scale\[5\] _0061_
+ sky130_fd_sc_hd__or3_1
X_0565_ VPWR VGND VGND VPWR _0123_ _0121_ _0122_ sky130_fd_sc_hd__or2_1
X_0634_ VPWR VGND _0189_ _0186_ _0166_ _0162_ net22 VGND VPWR sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_3_Right_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0617_ VGND VPWR _0171_ _0172_ net10 VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0548_ VPWR VGND VGND VPWR _0084_ _0107_ _0088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_76 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0882_ VPWR VGND VPWR VGND _0383_ _0423_ _0384_ _0381_ _0424_ sky130_fd_sc_hd__or4_1
X_0951_ VPWR VGND VGND VPWR _0471_ count\[22\] _0468_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0934_ VGND VPWR _0038_ _0458_ net13 _0459_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0865_ VPWR VGND VPWR VGND _0405_ _0062_ count\[7\] _0407_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_75 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0796_ VPWR VGND _0342_ net21 true_scale\[23\] VPWR VGND sky130_fd_sc_hd__and2_1
X_0581_ VPWR VGND VGND VPWR _0137_ _0136_ _0138_ sky130_fd_sc_hd__nand2b_1
X_0650_ VGND VPWR _0204_ _0191_ _0203_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0917_ VGND VPWR _0448_ count\[11\] count\[10\] _0444_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0848_ VPWR VGND true_scale\[12\] true_scale\[13\] _0064_ _0390_ true_scale\[14\]
+ VPWR VGND sky130_fd_sc_hd__o31ai_1
X_0779_ VPWR VGND VPWR VGND _0324_ true_scale\[22\] net21 _0017_ _0325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_54 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_98 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0633_ VPWR VGND VGND VPWR _0185_ _0188_ _0187_ sky130_fd_sc_hd__nand2_1
X_0702_ VPWR VGND VGND VPWR _0239_ _0242_ _0238_ _0253_ sky130_fd_sc_hd__o21a_1
X_0495_ VPWR VGND VPWR VGND _0060_ net10 sky130_fd_sc_hd__inv_6
X_0564_ VGND VPWR _0122_ _0103_ _0101_ _0120_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_0_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_59 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_17_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Right_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0616_ VPWR VGND VGND VPWR _0171_ _0169_ _0170_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0547_ VGND VPWR VPWR VGND _0092_ _0106_ _0104_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_31_Right_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Right_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_31_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_177 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_26_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0881_ VPWR VGND VPWR VGND _0389_ _0422_ _0392_ _0386_ _0423_ sky130_fd_sc_hd__or4_1
X_0950_ VPWR VGND VGND VPWR count\[22\] _0470_ _0468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_2_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0933_ VPWR VGND VGND VPWR _0459_ count\[16\] _0456_ sky130_fd_sc_hd__or2_1
X_0864_ VGND VPWR _0406_ _0062_ count\[7\] _0405_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0795_ VPWR VGND VGND VPWR _0336_ _0337_ _0341_ _0339_ sky130_fd_sc_hd__nand3_1
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0580_ VGND VPWR VGND VPWR _0118_ _0114_ _0119_ _0137_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0916_ VGND VPWR _0032_ _0446_ net14 _0447_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0847_ VGND VPWR _0388_ _0389_ count\[14\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0778_ _0325_ _0303_ _0312_ _0323_ net15 VPWR VGND VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_0_20_66 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0632_ VPWR VGND VPWR VGND _0166_ _0162_ _0186_ _0187_ sky130_fd_sc_hd__a21o_1
X_0563_ VPWR VGND VPWR VGND _0103_ _0101_ _0120_ _0121_ sky130_fd_sc_hd__a21oi_1
X_0701_ VPWR VGND VGND VPWR _0249_ _0251_ _0252_ sky130_fd_sc_hd__nor2_1
X_0494_ VPWR VGND VPWR VGND _0059_ net7 sky130_fd_sc_hd__inv_2
XFILLER_0_9_96 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_34_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0615_ VGND VPWR _0170_ net17 net7 net9 VPWR VGND sky130_fd_sc_hd__and3_1
X_0546_ VPWR VGND VGND VPWR _0092_ _0104_ _0105_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1029_ count\[26\] net26 _0048_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_31_189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_22_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0529_ net20 _0088_ net4 net18 VPWR VGND VPWR VGND sky130_fd_sc_hd__and3_2
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ VPWR VGND VPWR VGND _0397_ _0421_ _0399_ _0394_ _0422_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_37_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_18_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0932_ VPWR VGND VGND VPWR count\[16\] _0458_ _0456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0863_ VPWR VGND VGND VPWR true_scale\[8\] _0405_ _0061_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_21_Left_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0794_ VPWR VGND VPWR VGND _0339_ _0337_ _0336_ _0340_ sky130_fd_sc_hd__a21o_1
X_0915_ VPWR VGND VGND VPWR _0447_ count\[10\] _0444_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0846_ VPWR VGND VGND VPWR _0067_ _0387_ _0388_ sky130_fd_sc_hd__nor2_1
X_0777_ VGND VPWR _0312_ _0323_ _0324_ _0303_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_0700_ VPWR VGND VGND VPWR _0248_ _0235_ _0233_ _0251_ sky130_fd_sc_hd__nor3_1
X_0631_ VGND VPWR _0186_ _0158_ _0156_ _0184_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0562_ VGND VPWR _0119_ _0120_ _0114_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0493_ VPWR VGND VPWR VGND _0058_ net20 sky130_fd_sc_hd__inv_2
X_0829_ VGND VPWR _0370_ _0371_ count\[20\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_184 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_40_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0614_ VPWR VGND VPWR VGND net17 net7 net9 _0169_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_7_Right_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0545_ VGND VPWR _0102_ _0104_ _0084_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_1028_ count\[25\] net27 _0047_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0528_ VGND VPWR VPWR VGND _0004_ _0087_ net16 true_scale\[9\] sky130_fd_sc_hd__mux2_1
X_0931_ _0456_ _0457_ _0037_ net13 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0862_ VGND VPWR _0403_ _0404_ count\[8\] VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_219 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_23_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0793_ VPWR VGND _0339_ _0320_ _0300_ _0298_ _0338_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0914_ VPWR VGND VGND VPWR count\[10\] _0446_ _0444_ sky130_fd_sc_hd__nand2_1
X_0845_ VPWR VGND _0387_ _0066_ true_scale\[15\] VPWR VGND sky130_fd_sc_hd__and2_1
X_0776_ VPWR VGND VGND VPWR _0321_ _0322_ _0323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0630_ VPWR VGND VPWR VGND _0158_ _0156_ _0184_ _0185_ sky130_fd_sc_hd__a21o_1
X_0492_ VPWR VGND VPWR VGND _0057_ net19 sky130_fd_sc_hd__inv_2
X_0561_ VGND VPWR _0119_ _0116_ _0117_ VPWR VGND sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0828_ VGND VPWR VPWR VGND true_scale\[21\] _0370_ _0070_ sky130_fd_sc_hd__xor2_1
X_0759_ VGND VPWR VPWR VGND _0286_ _0267_ _0285_ _0307_ sky130_fd_sc_hd__or3b_1
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0613_ VPWR VGND _0008_ _0167_ _0166_ net16 _0168_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_25_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0544_ VPWR VGND VGND VPWR _0103_ _0085_ _0102_ sky130_fd_sc_hd__or2_1
X_1027_ count\[24\] net26 _0046_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0527_ VGND VPWR VPWR VGND _0087_ _0059_ _0082_ _0086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0930_ VPWR VGND VGND VPWR _0457_ count\[15\] _0454_ sky130_fd_sc_hd__or2_1
X_0861_ VGND VPWR VPWR VGND true_scale\[9\] _0403_ _0062_ sky130_fd_sc_hd__xor2_1
X_0792_ VPWR VGND VGND VPWR _0303_ _0322_ _0338_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_29_Right_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0913_ _0444_ _0445_ _0031_ net11 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0844_ VGND VPWR _0385_ _0386_ count\[15\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0775_ VPWR VGND VPWR VGND _0300_ _0298_ _0320_ _0322_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0560_ VPWR VGND VGND VPWR _0116_ _0117_ _0118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_78 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0491_ VPWR VGND VPWR VGND _0056_ net21 sky130_fd_sc_hd__inv_2
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_10_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0758_ VPWR VGND VPWR VGND _0186_ _0306_ _0225_ _0160_ _0185_ _0207_ sky130_fd_sc_hd__a2111o_1
X_0827_ VGND VPWR VPWR VGND count\[21\] _0369_ _0368_ sky130_fd_sc_hd__xor2_1
X_0689_ VPWR VGND VPWR VGND _0223_ _0206_ _0224_ _0241_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0612_ VPWR VGND _0168_ net22 true_scale\[13\] VPWR VGND sky130_fd_sc_hd__and2_1
X_0543_ VGND VPWR _0100_ _0102_ _0094_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_1026_ count\[23\] net29 _0045_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_167 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_30_181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_13_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0526_ VGND VPWR VGND VPWR net7 _0086_ net6 sky130_fd_sc_hd__xor2_4
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ count\[6\] net23 _0028_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0509_ VPWR VGND VPWR VGND _0074_ true_scale\[26\] _0073_ sky130_fd_sc_hd__or2_2
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0860_ VPWR VGND VPWR VGND _0400_ _0063_ count\[9\] _0402_ sky130_fd_sc_hd__a21oi_1
X_0791_ VGND VPWR VPWR VGND _0337_ _0323_ _0305_ _0308_ _0309_ _0310_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_14_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ true_scale\[13\] net24 _0008_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0912_ VPWR VGND VGND VPWR _0445_ count\[9\] _0442_ sky130_fd_sc_hd__or2_1
X_0843_ VGND VPWR _0067_ _0385_ true_scale\[16\] VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0774_ VGND VPWR _0321_ _0300_ _0298_ _0320_ VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0490_ VPWR VGND VPWR VGND _0055_ signal_clk_out sky130_fd_sc_hd__inv_2
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0688_ VGND VPWR VGND VPWR _0240_ _0187_ _0207_ _0185_ _0225_ sky130_fd_sc_hd__a211o_1
X_0826_ VPWR VGND VGND VPWR _0071_ _0368_ _0367_ sky130_fd_sc_hd__nand2_1
X_0757_ VPWR VGND VGND VPWR _0303_ _0304_ _0305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0611_ VGND VPWR _0161_ _0165_ _0167_ _0160_ VPWR VGND sky130_fd_sc_hd__o21ai_1
X_0542_ VPWR VGND VGND VPWR _0094_ _0101_ _0100_ sky130_fd_sc_hd__nand2_1
X_1025_ count\[22\] net29 _0044_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_28_Left_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_16_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_16_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0809_ VPWR VGND VGND VPWR _0060_ _0351_ net15 _0353_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_160 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_6_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0525_ VPWR VGND VGND VPWR net6 _0085_ net7 sky130_fd_sc_hd__nand2_1
X_1008_ count\[5\] net23 _0027_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_90 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_36_208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_12_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_79 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_41_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0508_ VGND VPWR VPWR VGND true_scale\[25\] _0072_ true_scale\[24\] _0073_ sky130_fd_sc_hd__or3_2
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_23_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0790_ VPWR VGND VGND VPWR _0334_ _0336_ _0335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_13_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ true_scale\[12\] net24 _0007_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0911_ _0444_ count\[9\] count\[7\] count\[8\] _0438_ VGND VPWR VPWR VGND sky130_fd_sc_hd__and4_1
X_0842_ VPWR VGND VPWR VGND _0382_ _0068_ count\[16\] _0384_ sky130_fd_sc_hd__a21oi_1
X_0773_ VGND VPWR VPWR VGND _0191_ _0320_ _0318_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_0825_ VGND VPWR _0070_ true_scale\[22\] _0367_ true_scale\[21\] VPWR VGND sky130_fd_sc_hd__o21ai_1
X_0756_ VPWR VGND _0304_ _0302_ _0301_ VPWR VGND sky130_fd_sc_hd__and2_1
X_0687_ VGND VPWR VPWR VGND _0236_ _0239_ _0237_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0610_ VGND VPWR VGND VPWR _0161_ _0160_ _0142_ _0163_ _0164_ _0166_ sky130_fd_sc_hd__a311o_1
X_0541_ VGND VPWR _0100_ _0096_ _0098_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_1024_ count\[21\] net26 _0043_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0808_ VGND VPWR VGND VPWR _0352_ _0343_ net10 _0351_ sky130_fd_sc_hd__a21bo_1
X_0739_ VPWR VGND VPWR VGND _0288_ _0287_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_206 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0524_ VPWR VGND _0084_ net7 net6 VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_0_6_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1007_ count\[4\] net23 _0026_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0507_ VPWR VGND VGND VPWR _0072_ true_scale\[23\] _0071_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ true_scale\[11\] net24 _0006_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_18_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_0772_ VPWR VGND VPWR VGND _0319_ _0318_ sky130_fd_sc_hd__inv_2
X_0910_ _0442_ _0443_ _0030_ net11 VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
X_0841_ VGND VPWR _0383_ _0068_ count\[16\] _0382_ VPWR VGND sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_25_Right_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_40_80 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0824_ VPWR VGND VPWR VGND _0364_ _0072_ count\[22\] _0366_ sky130_fd_sc_hd__a21oi_1
X_0755_ VPWR VGND VGND VPWR _0301_ _0302_ _0303_ sky130_fd_sc_hd__nor2_1
X_0686_ VPWR VGND VGND VPWR _0236_ _0237_ _0238_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_25_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0540_ VPWR VGND VGND VPWR _0099_ _0095_ _0098_ sky130_fd_sc_hd__or2_1
X_1023_ count\[20\] net26 _0042_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_0807_ VPWR VGND _0351_ _0346_ _0340_ _0334_ _0345_ VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_0_24_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0738_ VGND VPWR _0284_ _0287_ _0283_ VPWR VGND sky130_fd_sc_hd__xnor2_1
X_0669_ VPWR VGND _0222_ _0221_ _0211_ VPWR VGND sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_2_Right_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0523_ VGND VPWR VPWR VGND _0003_ _0083_ net16 true_scale\[8\] sky130_fd_sc_hd__mux2_1
X_1006_ count\[3\] net23 _0025_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0506_ VPWR VGND VPWR VGND true_scale\[22\] _0070_ true_scale\[21\] _0071_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_32_213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_32_224 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ true_scale\[10\] net24 _0005_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_240 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0771_ VPWR VGND VGND VPWR _0318_ _0316_ _0317_ sky130_fd_sc_hd__or2_1
X_0840_ VPWR VGND true_scale\[15\] true_scale\[16\] _0066_ _0382_ true_scale\[17\]
+ VPWR VGND sky130_fd_sc_hd__o31ai_1
XFILLER_0_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ VGND VPWR VGND VPWR _0050_ count\[28\] _0481_ _0482_ net12 sky130_fd_sc_hd__o211a_1
XFILLER_0_4_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_37_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0685_ VGND VPWR VGND VPWR _0237_ _0221_ _0211_ _0220_ sky130_fd_sc_hd__a21bo_1
X_0823_ VGND VPWR _0365_ _0072_ count\[22\] _0364_ VPWR VGND sky130_fd_sc_hd__and3_1
X_0754_ VPWR VGND VPWR VGND _0282_ _0147_ _0281_ _0302_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_19_135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_19_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1022_ count\[19\] net26 _0041_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_108 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_0668_ VGND VPWR _0221_ _0218_ _0219_ VPWR VGND sky130_fd_sc_hd__xnor2_2
X_0737_ VPWR VGND VGND VPWR _0283_ _0284_ _0286_ sky130_fd_sc_hd__nor2_1
X_0806_ VPWR VGND VGND VPWR true_scale\[24\] net15 _0350_ _0019_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0599_ VPWR VGND VPWR VGND _0135_ _0128_ _0134_ _0155_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0522_ VGND VPWR VPWR VGND net6 _0083_ _0082_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_16_Left_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_1005_ count\[2\] net23 _0024_ VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_35_211 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_35_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_26_200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_0505_ VPWR VGND VGND VPWR _0070_ true_scale\[20\] _0069_ sky130_fd_sc_hd__or2_1
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_26U9NK c1_n3146_n1500# m3_n3186_n1540#
X0 c1_n3146_n1500# m3_n3186_n1540# sky130_fd_pr__cap_mim_m3_1 l=15 w=30
.ends

.subckt sky130_fd_pr__pfet_01v8_AXJJQ9 a_158_n197# a_n874_n197# a_n416_n100# a_874_n100#
+ w_n968_n200# a_n358_n197# a_358_n100# a_416_n197# a_n100_n197# a_100_n100# a_n674_n100#
+ a_n158_n100# a_n616_n197# a_674_n197# a_616_n100# a_n932_n100#
X0 a_874_n100# a_674_n197# a_616_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1 a_n158_n100# a_n358_n197# a_n416_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 a_100_n100# a_n100_n197# a_n158_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3 a_n674_n100# a_n874_n197# a_n932_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X4 a_616_n100# a_416_n197# a_358_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X5 a_358_n100# a_158_n197# a_100_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X6 a_n416_n100# a_n616_n197# a_n674_n100# w_n968_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_HD5U9F a_n129_n150# a_n221_n150# a_63_n150# a_111_172#
+ a_n33_n150# a_n81_172# a_159_n150# a_15_n238# a_n177_n238# VSUBS
X0 a_159_n150# a_111_172# a_63_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.465 pd=3.62 as=0.2475 ps=1.83 w=1.5 l=0.15
X1 a_63_n150# a_15_n238# a_n33_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=0.15
X2 a_n129_n150# a_n177_n238# a_n221_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.465 ps=3.62 w=1.5 l=0.15
X3 a_n33_n150# a_n81_172# a_n129_n150# VSUBS sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_5VPKLS a_n29_n100# a_487_n100# a_n229_n188# a_287_n188#
+ a_n287_n100# a_n487_n188# a_229_n100# a_n545_n100# a_29_n188# VSUBS
X0 a_n287_n100# a_n487_n188# a_n545_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1 a_n29_n100# a_n229_n188# a_n287_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 a_229_n100# a_29_n188# a_n29_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3 a_487_n100# a_287_n188# a_229_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_99C25S a_n229_n1597# a_n545_n1500# a_n29_n1500# a_229_n1500#
+ a_287_n1597# a_29_n1597# a_n487_n1597# a_487_n1500# a_n287_n1500# w_n581_n1600#
X0 a_487_n1500# a_287_n1597# a_229_n1500# w_n581_n1600# sky130_fd_pr__pfet_01v8 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X1 a_n287_n1500# a_n487_n1597# a_n545_n1500# w_n581_n1600# sky130_fd_pr__pfet_01v8 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X2 a_n29_n1500# a_n229_n1597# a_n287_n1500# w_n581_n1600# sky130_fd_pr__pfet_01v8 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
X3 a_229_n1500# a_29_n1597# a_n29_n1500# w_n581_n1600# sky130_fd_pr__pfet_01v8 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_MMM6UU a_n287_n500# a_n487_n588# a_745_n500# a_545_n588#
+ a_229_n500# a_n545_n500# a_29_n588# a_n745_n588# a_n29_n500# a_487_n500# a_n229_n588#
+ a_287_n588# a_n803_n500# VSUBS
X0 a_487_n500# a_287_n588# a_229_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_745_n500# a_545_n588# a_487_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X2 a_n29_n500# a_n229_n588# a_n287_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_229_n500# a_29_n588# a_n29_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_n545_n500# a_n745_n588# a_n803_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X5 a_n287_n500# a_n487_n588# a_n545_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt buffer vd ib out in gnd
Xsky130_fd_pr__cap_mim_m3_1_26U9NK_0 out d sky130_fd_pr__cap_mim_m3_1_26U9NK
Xsky130_fd_pr__pfet_01v8_AXJJQ9_0 a vd a a vd a vd a a a vd vd a a a vd sky130_fd_pr__pfet_01v8_AXJJQ9
Xsky130_fd_pr__pfet_01v8_AXJJQ9_1 b b vd vd vd b b b b vd b b b vd vd b sky130_fd_pr__pfet_01v8_AXJJQ9
Xsky130_fd_pr__nfet_01v8_HD5U9F_1 a a b b c out b in a gnd sky130_fd_pr__nfet_01v8_HD5U9F
Xsky130_fd_pr__nfet_01v8_5VPKLS_0 gnd c ib c ib ib c ib ib gnd sky130_fd_pr__nfet_01v8_5VPKLS
Xsky130_fd_pr__pfet_01v8_99C25S_0 a d vd d d a d d d vd sky130_fd_pr__pfet_01v8_99C25S
Xsky130_fd_pr__pfet_01v8_99C25S_1 b out vd out out b out out out vd sky130_fd_pr__pfet_01v8_99C25S
XXM10 d d gnd gnd out gnd d gnd gnd gnd d d gnd gnd sky130_fd_pr__nfet_01v8_MMM6UU
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_XMXTTL a_546_450# a_n118_450# a_546_n882#
+ a_n450_450# a_n450_n882# a_n284_n882# a_n118_n882# a_n616_450# a_380_n882# a_48_450#
+ a_380_450# a_n616_n882# a_214_n882# a_214_450# a_n284_450# a_48_n882# VSUBS
X0 a_n616_450# a_n616_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.66
X1 a_380_450# a_380_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.66
X2 a_546_450# a_546_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.66
X3 a_214_450# a_214_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.66
X4 a_n284_450# a_n284_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.66
X5 a_n450_450# a_n450_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.66
X6 a_48_450# a_48_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.66
X7 a_n118_450# a_n118_n882# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=4.66
.ends

.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.2132 ps=1.67 w=1 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 VPWR a_1283_21# a_1847_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 Q_N a_1847_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_1283_21# a_1847_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X13 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X17 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X18 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X19 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X20 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2132 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X26 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X27 Q_N a_1847_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X28 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X29 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_XGSNAL a_n33_n397# a_n73_n300# a_15_n300# w_n211_n519#
X0 a_15_n300# a_n33_n397# a_n73_n300# w_n211_n519# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_QABHPF a_546_200# a_n118_200# a_546_n632#
+ a_n450_200# a_n450_n632# a_n284_n632# a_n118_n632# a_n616_200# a_48_200# a_380_n632#
+ a_380_200# a_n616_n632# a_214_n632# a_214_200# a_n284_200# a_48_n632# VSUBS
X0 a_48_200# a_48_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2.16
X1 a_n450_200# a_n450_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2.16
X2 a_n118_200# a_n118_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2.16
X3 a_n616_200# a_n616_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2.16
X4 a_380_200# a_380_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2.16
X5 a_546_200# a_546_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2.16
X6 a_214_200# a_214_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2.16
X7 a_n284_200# a_n284_n632# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=2.16
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_A4KLY5 c1_n2866_n2720# m3_n2906_n2760#
X0 c1_n2866_n2720# m3_n2906_n2760# sky130_fd_pr__cap_mim_m3_1 l=27.2 w=27.2
.ends

.subckt sigma-delta out vpwr clk reset_b_dff gnd vd in
Xsky130_fd_pr__res_xhigh_po_0p35_XMXTTL_1 m1_n1920_4820# m1_n2580_4820# in_int m1_n2940_4820#
+ m1_n2760_3480# m1_n2760_3480# m1_n2420_3480# m1_n2940_4820# m1_n2100_3480# m1_n2260_4820#
+ m1_n1920_4820# in m1_n2100_3480# m1_n2260_4820# m1_n2580_4820# m1_n2420_3480# gnd
+ sky130_fd_pr__res_xhigh_po_0p35_XMXTTL
Xx1 clk x1/D reset_b_dff gnd gnd vpwr vpwr x1/Q out sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_pr__res_xhigh_po_0p35_XMXTTL_2 m1_n440_4820# m1_n1100_4820# x1/Q m1_n1440_4820#
+ m1_n1260_3480# m1_n1260_3480# m1_n940_3480# m1_n1440_4820# m1_n620_3480# m1_n780_4820#
+ m1_n440_4820# in_int m1_n620_3480# m1_n780_4820# m1_n1100_4820# m1_n940_3480# gnd
+ sky130_fd_pr__res_xhigh_po_0p35_XMXTTL
Xsky130_fd_pr__nfet_01v8_648S5X_0 x1/D in_comp gnd gnd sky130_fd_pr__nfet_01v8_648S5X
XXP1 in_comp x1/D vd vd sky130_fd_pr__pfet_01v8_XGSNAL
Xsky130_fd_pr__res_xhigh_po_0p35_QABHPF_0 in_comp m1_n2360_2660# m1_n1860_1820# m1_n2700_2660#
+ m1_n2860_1820# m1_n2520_1820# m1_n2520_1820# in_int m1_n2360_2660# m1_n1860_1820#
+ m1_n2040_2660# m1_n2860_1820# m1_n2200_1820# m1_n2040_2660# m1_n2700_2660# m1_n2200_1820#
+ gnd sky130_fd_pr__res_xhigh_po_0p35_QABHPF
Xsky130_fd_pr__cap_mim_m3_1_A4KLY5_0 in_comp gnd sky130_fd_pr__cap_mim_m3_1_A4KLY5
Xsky130_fd_pr__cap_mim_m3_1_A4KLY5_1 in_int gnd sky130_fd_pr__cap_mim_m3_1_A4KLY5
.ends

.subckt tt_um_hugodiasg_temp_sensor_clock_divider clk ena rst_n ua[0] ua[1] ua[2]
+ ua[3] ua[4] ua[5] ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5]
+ ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6]
+ uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6]
+ uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6]
+ uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] VDPWR VGND
Xsensor_0 VDPWR ua[3] sensor_0/vtd VGND sensor
Xclock_divider_0 clk uo_out[0] rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4]
+ ui_in[5] ui_in[6] ui_in[7] VDPWR VGND clock_divider
Xbuffer_0 VDPWR ua[2] ua[1] ua[3] VGND buffer
Xsigma-delta_0 uo_out[7] VDPWR clk VDPWR VGND VDPWR ua[0] sigma-delta
.ends

